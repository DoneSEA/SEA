`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gewdhL/w1TouB0JjuZHJxluLgazZ0MDhwTiI0DySlF2H3xd6FRSfzLr57O3qUZ5eGvZn9G1HUOcz
yxVE1Ft6ug==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kNkvEiBddZ56G5aF+XS7ob2Nhv2j+6nmCRkSoQq0oirSRWu0r3CeEeHNjMTnlz141inTsI0Z6BWi
mSQVN+vnta1jke0Bk4Stt+1AehqmzqWBhIHNifuASwGS7djtqVZP4SiTYyIWLtw2ytc2NIoTTIPD
p8KuPz5sCnz/rVbTGrU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PQCKWrqcONejuC35aWg8w9DioCraSLD3jpWb1GhpUCgcaZ0iGFYF6zyTQ9UbFoUruOqUsK4NCVSk
hplF/dXRzE4vE39sCsuYrnlvsXoMvw5omH6qSVsPw0ouHfl9A2UJZkAWOT/cmxzDUB2Nwx6oDebh
LR1vONCseE7uyR5RxjiK0JeDjP0hoBNJoC8RfEDbHpmrb9nOAmibt1Ub/3ax1qZCSXM9KLwO8O6m
3xVW+RxfWvYY4vl1SaNWMWCqoW8nl6bPZ2E3eaXRj1MmReX5VOJjdR+D+uJyoaWNDJWHitCvsaop
vIHRQS6GhW6gQDoyFrOee9vd8Mk5vO4zHSkoCQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EnheuADwC+rXRbRg9Il4ySLQns8VKTnppIVWIV7/j1q3n5T9ImVRYukn1hvdbcKoYxtL+2UcCg96
5OeU5Cmw2OktWg+nXUEQsGpMI/HtDbo51bYU08HKrrfZfLFzJht2bJQKefep8XtA+PBarinw89ic
y5pRbW5e+RK1wq2fpuZ/aad4nPvIc4RQLnDGpE3/KsO8mmLVobPkafsCgRcjsOloyEh2SIKI0L3S
bM1yoTNj3PBKHQ+Fg5c57g4tgtPWlOZoENX18yDgBTaLFQz2pRFtbb1TFYKxNIWOk5nYHwQhWhGV
7FfMa5zdnsgLXGK6/E4ssQcSyIcY1ZJqqeKUWw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
w+as5hQm6N6F6rMbvXzBeWbsgKQk/heHkIxjXuTz4RzbjzgbTltcE8Flz3fkoKf5N7ML5dxsjo9D
ssHdLG4rf7XR8V4jTftZ++etToKtPnQBCB9DKi1yN533S5ArNcUfnE3UNrkiVdemu8VNDcPhkNGG
T6L1X+PWyuW9l0Qj2VQM4rosaZCg7fijmq6q9IbXnhPGGcvP+YH+yhPpUX2y8PH6GVZMCdpdUpkd
gEm8oLFSJ28Q7zZvqQZsrdEIlThY2i1c8NDuhS8NDtOmlumPhbPr7rKYBAwl6DCIXO+CqE2a8X/c
qpIBWTRvLyaD7BcA7XDCyMfCZy/mq8fZ6rIrOQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ebIGhwOoK6b2Regd2ZidBmefLC1qWrjb2ixldIHZBv9r8mN994nK0bA5i2yPW5FfOgPszrabIv2T
d9dzSTELNwamhC6udZmN9sBwlaEVqro7zC0hwc9PBph7uwSv+FXYBFkXpe9DnpJTZbUvUeThstgk
RdebU+EnQryZ0UpzZ2A=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XnwajLd9gtUhj/hQ3dArVFrFrrTuWhrvu+kPxwrOfm2NgABPJQFBXwBwCw2jjlhA7jCVcZI4CRq8
GHr5uL3LcoFEL49z34pdL9z8W+zlAFZZl/rnslm3zKW6HpX5Z9zjmS0PThKZoMBpBHWSEKjmXjSE
t+thGVHHTSqS9h2Uo8qpx2g2fY7ITBA2F2G3aajNf+o5hHTA5QnC/87hlfZzNl7Redk6aQRYCgB8
LIJBeO59sYe3aKg/vswdYeXiRdd8b45eVOvTT4iKpa1ExnseAad7tGfp2qVyT4QrHVx9jSYd05Mu
8Dlg+1UQcbk2h4Q0cJ7WGdpp1ljWsx8j2GPrQw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
Kueiqp3scnBkX5wNz6pkll+oz4mC9E58OJXFNScWRYtCzd8FwcTT5wwnYIoOWyO3SMHOd1NFN78z
GyvS2+mYl9XObeNn2dCWfhZ78N+lnWAQYNDcdsdHupvvPD+OcrDa/Cmvdnvzo+YcWXKEEfoDnW/T
7L+cEgmwwOgfH2QI0bjovCU/2xsdHqsr1yqSV1ODn8YiJgtvd/kJ8gtEVHdrcupxdYQKY/h9woP0
KiZGO0ptkI5r4UEvPLowYYnWEzIJ7jXK5qYJUd87HiiB6Qc+esT/bakKYLo5CPj4bl/otlzZZ0hz
p8Uaat3cpmP/WoRL6Hjmex8YhGS/CKi/YA+OG/dK789WUL4Oynu8iRxz6QcUioe6JW4wSlSKbrKu
NB3BdwBsqIRC/tJx+elWTkpjZYbKgGR9LuHe6yPhcoev58aBvvcYnayYuRUvmVD3ZIKRe3kO9oWg
St7XbdZjmyvgs3S7sU5Ph5TCrtjJHQo6dcGE/hjxodbEIizEo9JrJXhvFpPbuCxQpNaxFtIid4jM
To4rM2aZd7xKdC/Nd/JndAmDBs+u2SYceAkmLKFA8h6Dv7X3hNkOymxCVOez6y4rQRM8ZR/ahxAs
6o9pi294v/3ZFrJm0kUd/BGujs/8R+N2U9q8ivm4b9wMAZ8oHbknJ2j2cGkAV1whSypj9EGyAGyl
Uj7++mTELI487AOCs8/qbeaGC2DjA5ErLqGCVDNuuIB9mvSCoBQDCjMuIq589mga9Nu2xz5poKO0
kW7IbK00cRUt7gf0dbIW57y8+6O/6jEVAiAeySknD9tQ//Ro0j9A3ZOqFwhagfrOasD978i4z2BG
rqnRfZnw3HQn3zdiQioTViHnO+1pL3WKMmFRGtX73XDc/MtYGo4y9oXPzTsn7WGRsaUmyIMauRz0
MtnhRUDVgDRt2+olPvcl2VZ2yADiC7v8yZTWkEg6W3LZTB5huwR7/W4M2PUiFThmfSNCMjkhgKOD
u8yeCfClTi+lMlC9yCI6Rg5NldOra1ot48mWc9ZOcpVALa1VwZ7WRrSzUUI4P1cIJeX/Hu4wZNFe
OPPNiIVDThHODXWaLqpih6RF+NRBxT9wTy0OsGDhAqrY9Ho695c5EBoGlPIleRr8k8YBZUx0IK41
GoZOAPIB/Uu6tqsaQgoC65f6euPzSy7lrMVihpmQBqXZwb25pc+vadOEr25PRYs/6QvXp+c+sDqs
fv2FtvLO0Gmt5lnpp5FkaHaMvSTk3tubNJEA7qU7MISPOT88FnXMw7p0EiV5SvvgizsXzWY7uPoa
HyqqZNPrAcz4RIvee0QDuIohWOEiaowfqerYzRLGJD6Up45oCe+3yblW5fnkUgoueAjN58Zd2Wcr
udcQmnmuD57FvREw4PIBzTrS+OBew6AGa7FgsEDnW/ATc6pCmIL+vGwvmc1RAq8fHMn3GhyGX7P7
6gQ6X0mUOaRzwLSJjiXytKfDbTUEwyEUaF1EODOhkNFXHtWT2p5Uui80d0sv65jOy4gVyizJ5xCL
AkGbglXVHVOj9zqQg+xOwm2ZzWLhM8opi3SZIUpGxomxt3GzM59O1sNUQFLBg+paZx2zLVob9qEM
drVLlg/Cly6uDKk+md4fIppRPNhTIQs/rO+JMMTsT2rkCfrouz6VQKIThKedfDf5cVU6InBDMYmM
/mNnvrmqhABqeCJP8tW8/o4F+S6VvX+euzr6qTeVlR6LfW4mSJD+qh8Qo7dACTPiRGmVxVd+LVmZ
uDrTFccJKrZCtjxfu4Ow+Co0MRgr+WN4AhZxgE6uz8NlT6hjadO+HybZo3ytisD5kDxVK6/hJMZi
fdCTyK+U/BcKFygalEzhvXTenWWOfxF6+oz0tpVBsJQOZHB2mFBMeSReQPXO/X1Zr8PHJBmvYfEd
vrptL3gShUJIwCc9agRuNXqOeD2gL3ru2qmgnU5pIO45CXkzKszzLJphuhs/RHwPBRK7bN8AFMBa
4p6BFukuDx61keUl+qUbzzoTARJuMatVXBhKXaDnFWbP2/dZkpYowxFbGXRxEm3FBRXl4DuRR2Zl
hm7qnXkis8fpyDmGAR+GvbkUtw3jB7WZCImL3DMVoUZ4Vju0e0zLyMvmQ5mUBqGWhGecufPkdJU2
YO3qPGJVEAovor1PTu4FOTNzLI1EFehUnaStNN6YaBYn8CwJH9uuT4O8xAbjY+rVxFd6oOByppPL
CBfTXVaMqS3Pi2+hJBwHYU57CSNCXBUS3Z4kx7z9Kl+FAtRGr8a+BcZUUeYk7y9QzXVwjbnEnLMs
/x6/b+F8IA32C7qB55zTUi8hwy/a5iz2gzibfXpZTj5Z2cZnvrzrLfW0qid4P4dHbGtROWCR93cC
BS1vnW9fIzt6jgYBLk5vt6YVC/RwArTJPxN41tGT19CJWlQkcCC+J0n9k4sf7T2iIJ+8aCKZZX08
q++05+FYgzLnMOrLHCq7wpDVomVtDlVO+5NuZIWJqs7UmkJmrc1XvUAdX7cBbkJK8TWH67HeOfsU
uf2TFmIU+7cG0VWgOi9JF7Rg7QHhvXHFgskJG32VkZH/+ivU+h3DQ7uoeS3vd3lxKRUPGkRRRsX+
KbYqB/usX/rMf+a/UFAT/SAmQ/o5755lz3keg+gVxOuN+Rnz17ZTZp4sR7PgfDc9NT4qkLSUKgR5
FqMX38Z8dQul6sA1sEwJBgRqQ/7+90deBTRy0hutW4p61JGdd+zTA8U9kdliywNeufnQQwi9bdkH
y9msW58Y/1u/YdCNXsRBZk4sa59509gpgHYPhMEt77d1xfT1xz+L2S2TQkOn6B/unn41hoCiv/Ej
/eZmwLMWD+RQp/Ekj3Dddgrd3ayuG+0xYRl+4k/PxyPxeimRwF3A8fxGw/WXeupbmw0q0fAJipDw
Pqgk+DdR/Gdrd1eLus3GkesyLtwGPBk2na5oBIeQ8TAoC4jEiVaLJNEC+3K1mptXClWN0n9h8hI+
10BUxOrPH8TlmG4m1uo+/Ng8JMTuMCGDYTISo3qIh3hLjftBiG7Gwn228vTsYUAIpbyMAMy6UaiL
tRJabdE6RD2uGT+a32c7cw3Q0AlA417VcPSqAPMbRMY0lSKLFcoC5EbKDupLOTA+sTgQa5vOJXYs
fJ1ducrd10ih6EpatTfzjb56NZPk93mBNjD0I5X7oxdkEY+gB8JCORW87BhqGZVqEmLDBte864sf
G7K9DwUlZqoyQH6BZHM1P1MMZCyoeHPY3+Vg0eKBOfa8GFuE2lMnsA3mPrlpQdFwN5puX9dK3yf7
GhIDjiIuwGxl2BKxYebOcJgWTNEjyPQ5xEcsvF1llhuUdLpwROpUOhX2Kv8//JN1bmVqi2HL3Y54
yT76LwCTjYvxG52ZUWXOoZlGe4+lAidUHtr+gcAcUkjMwuxH5BoLTTP4FJ3z38GxFecS3rs9JbY3
jqLrn5mUlvbBsFJsHbAZQbuCnermOkIy/lSjGJftJGe8AqNcUTCAxtoDn+PYD8f03jQeXiJ6M/iY
/CY3npnTBFW7iBfLDqh6P2UMSdW2XGDocLs8U5OaJlpZ2ccowNf+YUONiOFWOoG1/h3Iu1kTJQTK
wypCLWxbPdZPEGzSnYwutHCp+F9cezdvsNIedtzF53d25I+/pNoucsiiCKAsSgGrq/4dW0Tk6cSr
0hKLctbl59hDATL5bwe1uYJhwlfQB7vy/wz1StMOpe1KSk1JJb7p5LroPXir1SbB1goHkez1ZNaJ
sd1HivlsmZiNkbqHIuLSHjrQn+rnL/NVhxaP4GOq4x2nKHQeELVdq0KbgLx2zwd2qDfrwIJrl9M3
MGsi8vV65suSxyEEFq/qC4/l8GlPvmy67RCxxLypZALjXV2boQE+tjiqfC/Fo5QwCDvzeufQNmBc
TeaTQTYL05D3loZm7wZX+2CuRI380jvjFrdIh9SE9KxKC91pyFnBLzrgsBJ7MW3jurWzXOvfaMCQ
SZ6luDcC49RJXIspcE/BF4u4jH9Twf76aiPT6mUQhCjXGm58K8Nge+WzhPChiP1+VJcun8TbxZMI
rDnUaWZrXk5jTPoExaq6gzyxK25VBcZa8XhHa2+L/n5KL+3GbTgeQl+PyVPIavnwDCyqvaxJ1idp
7hdXlbCgtDfIWrWotaHTj0i7SiPsIZiboyGt9BQnPOUOUSosHQyiniFgQ5WUYLIYpilaEegd/dYr
iiWTzPR3qx6Z91u/5EPh+u960a9DSEOJIQ6+0PXXg1yjVvTbCsHP7RlpnFsdwAUfl5VOsyt3Cuvi
Evi4n7+zwIB8lUOwjnf8OEqWdy+15XKd/V84HL+QqVlIIdA60TmgSlvJTBAUhwM1BMT9hYwv4n5+
g7PQs8KiUoIgRYoUZ185m440Ex2378wbmmQ78dH0UN6mjSUjTM2MgpIk13wSy6cC5kT0i/gzE5AL
z2U0BcBtYbonGPi1JCgE5GlIxCK1bkbqY0eTZNCvnohYPU/g6jyhj8cba+AhnPCMTaGqkZlvC+qN
tlx1dHgrSCg9jXvDJJykZ3E7mDge4D13OSLWHkG2BCEkUuyzFwgQcB4gBIj5JfkCfeBzrcSZussc
tS6qiFX3+5I+4GYtOfgGHIdwANU67OvIMUdbB9N7OEUrLGK5I6LACWw+kNW4I52dIlRRI19zia2/
1CbwWcUgFTuinYa03U11b/XjNWkkpbUh0NDD+sMb3G++ucSfUwm6TIcpnV6p+LdcYz1prHVKeWBj
V+AB7MPLwm4pzIp4A6cwheOuE3VOxqlPJgCVE7LGSTaT4vsWKwjGAse16Rfs8dg1CfrSRhE1Lceo
KUWGscomxfG9FxkxacbBU13kzsTAgIF1RaWI4exe4fidGGAMnhz9nmQsT6NDUf8icAYOkBLKChn2
HWvuCdiINff+z3ninr0CCQjwY9EPSDNIbpIIFrIj40TZc4InvVRrHIoSFqEKRkPr+E+IlwH+REQK
SUOfEf984cE1MY5RoqINANzR8oOE5I+bbpZhKHwcZSfMEHEzm8fe56IEX20uJGshMhLTwttZwl6v
a6JN54S7/hl+uMGOS0KbqQQ4wQdIu3V0HNdg4vlyhO9JdTWgVqa/t0sBE5ecSYk0sZTQXJjMCHzW
X6/xQfNYmCu3kqEeF4UNJ2OkpuKZJ1EnykQqAk2/UVhwtKHWr5oEDHT20duTrijr0KNduEpUykzo
fv4OTdkxz4pUyR8DxcVAO0N+bWuQ07FGnFedkc7mTzZbLTn5D4pigTJC22hivA0QhGp2Xy1VyVek
vViZc0nIVB/R6gMQJ7ylm2CYs/7rKO13SmStIUGOYJdIfwMsa3gOyn/Z0aJfmG1+lG/dWslNWOPO
AYg2PjlWgCVLFauGx1h+FaxmgKeUvjv1KvMX+iwDNpOksi442ZQ9uOqUZs4gxSOc8moHObi1PtBf
3pbk+g3WzuczK3/28xiHf1Zdl6DXvvB29BOgtxOhD58h8mk42k9JaKDlnkM8of4XcuWWnqWldpa1
DLWbuOSalPg16AUbSqpbWcKD5Z0NFSZ51N5CyWkjCOmSVydCChx1g+IWDTB6FVg9fgVAV1nMuHYf
m9OEGd7ZLkTPe42aaqKfuOBDoNYPwBcWwxpWpgchndSkEpgwmfDWpGDH9LpBlhWFiRHdRIDCvlbh
o54SuoWUTJDsrsQPOEguWil5/6Dm43Z6XyEKF1arLg3fw+I2Y9PmJVyninscnGVCdeh/fi4MsRYW
XndT7IKnrDgWi4VafWSI4zuk9+xIO95OOgutM5uwOApsJoj2edGQzqn6Co/VLlxSUVJnU04n84Rg
EymyxpnEJ5uG4kIU89SomB3vtUF3qkghvBaiqAJF5kIq9N3YVggf2/yoiyHUDmblXr+Le3YBIV4o
F1j2jSRPKYHZLcBbcEGnlt1KAgb8nRmTNkTNw1ZCNYrDtYcgrbZ6YHXNJCce0+7pYZzM5HAPaaz+
FXLU2MIHFpn45pyEQkRUltZv//ZcmHweiaVmzrrpy8zg+uOPEltBTN+Gmnq0a2/SBRhmieXF79ri
zujGqvn7zZuOTvVG2CB7YjDPhWxAgoNetHQybgSXpUk9TJeICRN6w5si2Vf7R4DoW5KapOKtX1UE
xVFK87dpmQvgSrx6Ivyo9mVvK1EHI/yh2TcVpXf8tu62KbjCNaxOrTyZoIoWjXaS5lMC3O+JLtxb
JNUQN3a7AndVasfvXwD7+Y1jgcM+Q984dOotPblBDXSHNjjePH8vQjKfiPutlG3NuspfKzP4p+/Z
RESUogGFiNKN5Q5fUCzOi7OijTZsFCIHMgaHw1qHkfOVK4xdwnX8M5GV8Lvw7YWXyN990Yj8fV8g
sYysj/y07nyX8HUbZkEeojrRA/7dRrv9xbA/GD7jWhnrig4nK3RJfkfsZevBsqJ4703Q08qEcztZ
ojQSw3xM8kT1Uawi3XRpomfVNAXA5SPbBfPrNDqbUO8sBbakQe9a3oGebCbL1tPav2Pai2BJ1zmC
Au0f8vJrfSnXgzvOBcGZsyxyw8w2hOM9759ne6th+nP30s8DDIiDro+n5pKmzEV3ib9QGCXe2sRc
57rw4I4F//9k5/PIdXRsySV6gR9ug48/zU/oGZStMtSy3KkI/FrCkYtDsWvoC3MvKkyDrG6wm8DP
xx5Whl+9DCwsfSA3s8xvDwGnZxttQef9y6v5Xg10gwHEnMPuNWJvHB2Q71g1SL9kv/Ey9+MKM2rH
iMpDocdl680xhyFGkCgmYmUBRuOVfc3bRxadCPcqIJJrjm16m5i2/dJCQuUnKaKFoblUFYIvv9Rq
KCno1G5Lzkt/WHr+Ilxj3e+RohcK3OgkekPyljVIZlV/NC6AUxYhDJX7tZvXKKMtH2UbUOy+0YPx
2mJ/5dUiXwos6OmoygCPlaEfADW/6KdiO4YoYvNAy1KNWwZOZEfVajFdByn9EcT9W7DssRxYpE1D
wp0an5VUc0983hdLGydr/1fWjxcsHeBxEvuKz74izEcGswOawiKDm2zP9uUcRkP94wZjRsSvNpGD
8sH6AaZJe8hYW3EPuz+31WyCeTveafeiBgFx/jkH3nIGePzGieqy58Km/NwLqd2ltguurIXLRiuv
WeOTQ4/wuOa1ffmF/s022iF40DUJ86ByHZfhx6pHtUBTmesgiildjCXK8aZWaVOmvpe0/TDAzzRX
EK8XYDIc8jVJIIrCzeFPoSRPma0qP5Og6GnaBix9dUjC/exP9iE8XOJeCTotM9wcmQZocKvVISms
GhdMyAelC+e16Gz+3OS1phcH2NZZVLRsrgD3jiGf9GKIwZXYz+rYbnqU1EC5N+j9RR4EnrLUGncE
JflvsHS3CJ15HiqWhz9PIv/9c8LssuDABrR1Vcj8dSBpAgSr9EDK2zKGQvSkRSFHjSaTHh+qv/I9
yR0HNE/2X0zjRp2FfrEio7z0ktO/45AOL7PWLg6IvzE01ZCHSfDx4S70JzkBaDSIMB0tU2tgSTAB
/U0sHKRc5OSDnrsGaVYfsUCD1rvMTbO8VaAe5EW9jjtwr5A6aYlfPV2UEMokGK8Gz73zxLx42aIW
2Ch1ACqAIhHqRut/1m4q2Iu3JZmz85jA22ie7tbb+5eDH5HD8o7CWEN1wQP+9Qq1znslA/7wyFjI
bxvY+wp412bM/GNrRJLvTuIOc4TiX3I2q9W8ixgiBOCzo7sbiuJ9r82xLLUWeLfAr9vGUmGEP9tm
9OkBE8zsA3eXBXNwr6vOuqu9b0QC5jf5c+Lzf9HnTHFswpAULb1a9AZTZmJ3QYOTvXyh3iZ8ZVFJ
RagbGBE1GlSZntQhzXnY1Vr722h/tm1veku/I7O7GMJMFIPiwXGjLk64ugUdQ+0n99f5r4v4LSIl
wIWUSKCi1TMobWjgWNXp0YJrjtrJColjYTMY/i1eoKs6lVDsWAbg3yr6JbKzOwxEASDb+tybGtd7
g84WED4d20sIfahJPLGNmYthi/3r5kajq7lGncq6eCRRiHkFelptrBuBtW2z8TmGQIk7mERJdJYA
Hii0VapS7n10z0wtcynJSn2H9M2hMp6HiVZhqqMmB4vykcKCciHCQQTJaLbg/gw+PzuG+NbjJPTC
zgCw47IwAXdDZFOgiT6q5CKYBp3BxngTbGkTiSBEJS36ixMYB5R0c41g2RUHyCX7nCPvvLtp49q0
8XlcrHrvHRPGjff/B78zbudS5DI6InVPEDooF9YDeJcaIECPPI/NWlTZs1NsfR7xk3rDnF8W441Q
niKcbFSYfUIdHL0F5Dg7N/BP+RrI1Gq1FDSVleE0yTul+XyTJtUqZNnQ2xLIPXHpNR+xsRCsLr0w
xfcvyHSP/blVeg+xy7rt/AkUvhacjgCK/aP4R8TtUylaV19kG1ludg4cmTakvwJXcbwcCG6XQixK
LkSA/4H+4qbKb66BkHzXjP4+Y27eHOYJ3fnuRwqPG0Nt3ezanpXjhpvxtl31vDstVqufy9xTxvP6
fTeJqNO96bEqC22xToSLYgfUE7ZaT5FD3izPvgmQgsC3OGmV62cfraTvpiEEZwZ8pnn+HbkRnvAe
pFLJTrFZlepXN7WoSeR2M4plYOVh4WpBgxzJZLN9AAZlBQPUGTioD73LLD12nqZf0covQroj3pTd
TjC1MJOxVbfJy2P+2dBlUXTtRYN5lRSRRBoQb0pk9QduXXUkk3VJuFj9fb7mzTgtSas4DtP/CfR9
kmJ4BfHP0+1DfwK3hVFzvCitO/4mjvUbhlKCGJhbl43h3eGyhKYVFdwtjulUMuS05G4rMxFuHl+Q
pyjzGUo2BXNv9XhjuCI+cfa89yv/1cLuodsWWWMvBqqJI8Q/KCFUc8hsFOSyIu2CNaJ5WBobKhfr
sVILYJbViLcAuVAKVHNfSLnceOBV0PfGy5A67gNk+nDdD9c+FQMHB/lYj4wByjpl8EIrxBDVaOvp
Rdl1cJWLpGXLJVB/3ffdFwOfHF0rwMjQ0V1D71SqtKUT0d/Tdyj8KzZ3wWANjppExLQW1vHz36aD
M0rPC1TvhkWuECQ4s8Br2gEBvATzZVCOKYp0IO4KQhotEDJXFwxQ6iw/60Rnc3nxZGrys+FxAQ4t
90UmAdi5bGIkPf9xFydBaHvvzKdJTXO4bqbNzv8X2INdCWRMyr7i77rNDAll8wWjvOHgs9ZJ1jlh
qxq1aIwtUh379k70f9/aF6EeiKco3T6/vB4R1TvLG3OCdbanWkmq74rVfG1vShVVSKHz5a/e4yGd
x++kQ+A1xFYgH2P285fTga5SsJpnm+aZUWa6HfaquyccWsVubRPEXxKV1kh8ljhFWFflw0tRbDoX
L+qAXzZA2F3h10WdnjfxdH1fXthoZuyDegSd+0COk8ghO8zVltXeI+JuvOuT66WdHnYYlNH8xg7C
vp4WCmErMncBxw0bT6Q0HIwc9QILXOVmOqBjpH8FqoAOhwhxrQSLuZxHykpxwGlz4f2QM76whN0x
XF5kY5MGRHQ8u/zSP5eGuM21YkTTtUkSrVa9vdPg6SS9Q4QvkVi2qkmQONcKU6YeNrNJ6qpHEH8i
muupDvDA7r4GUOBcLYxkH91ebPWQBFWkLOO31R7Bilnj+ngfywK6Eh7YeTtGqq8Ku6At7WE9h++Q
Wip2Ip1gub1I7FEFxtlpRFa1dezlPlfwq4qPBxBuSLmeMmRXK2/oqAnckFRM8Qi0bL+Qe0tuksgC
E9JxpISeBrsO77j+syVTbwtebyyREutUinyCfDtncL8XX7d64pekX+wJY8DwjSyvYDtY4HlEsVl9
dfwdgBzIb8BBza2l81szRV9ABdmCQRkMIUdkiOpTiR7JeRDaJN0G9G082Q0UeTm9lsxumX3qL8gb
9oe4sBQkQ/HSO+cMG2MmCc0JKLwo2JKrNs0XyPTs79CSMqiXtTpInElM48meKbYWsAZSHj/mZeG1
PBIqfDPkMZ2x6AWN/7McxOJCN2ia75qdJV9DJesJWql6TIWeWwtAwyxG4Nwidi6EPaoVWYBMUxLY
XFLlDWIAraH8OvkfNciZ0it6gO8CJlJjAJ5XkbzgDToGilDXVO+dSW3Iwyorh0rzQw7OUlF/sgni
SuJs/LF0UJ3jiDA7UybfFahBA9algb4/e+6wyy6nG/2You/DCO0UeWcTvpb4C9f+VjSByjd/mmFN
CGVZ2GZ8860MJX+OIyTeCNzJjV0sUWYzv/8dyOWkiXd3ujBJp0Ux8gGQG4vqiBSqEfFuaGlEBD2e
b2V6Q0weP/rvT43dA+ISJXH+732CyiwXoaWVLg8DxzAGo2cSxXnsDrJvLV0oGLZvWmzmPygOgCUc
H7sl+1TSrJDo6zT+sVmwQUpSLqo2DhBv2mSBGfzVbPYX1ZkMOEkM2BVjZcNa7sWyRuDJ/SL7eRYn
ewvUmu5UadbNcFQCD7bf/w6MzluElBUR4RXfbOGT2sFoONHcglnqqLfSXSn69bwcZWV/4Nhk2cNq
CIGnyF76VKubZ9vRlNvW1QtJkw39AV2rsIH7qm/noxdDY2AIWbQzAEX0Q0v+C6LETfQPaJC5QbQV
qlHUqXVehnuzUWVAh2ush6h6m2gTFAmNxAQhakJ8xqIJpXuN7KIz2oMsm9jshzvNUuGY8399I+mj
VOjx7aq+RKTGRaB9TcMx1sJLw5HfU18NiRCG7l2wfWayDM281ESFSRNTdtFw8kqPDMryF8zn2Qz8
10k9rPy/kd1Kz4uo93L4leXTpW8XWI7TRpcGqy6kcbUJlm1U8fZ20R1UYiRe7SxFIjwzm9TbIPXr
DmS7+QJnG0rdzb9KH9epmrLfx8efnEP9lcstLwut53wKBoHuQgwMqqjxFbl6KWuYDqiysRXXUVvR
JXwk2T/o3N/WuDc+OlLbqOdjw7dilgI30ClvHo/QaJoTv0ZKz8jVJ7v0PK/xiV4Q3YIuBXPiDAfg
dJNHdRNoAjT4k8XFPvjzIOIpgggPY2COplU5eTXzwRiTWZpU+t2i7SA1md6LgfjO1LCZlcAmTNHv
Z/gnyl2AGBkm6AeMUBef9oZSiVxzCwJC9o4ggMVtijpz0FsqNoqeUPsQ7wOI3iBEnbvrQYZKRU5v
vu/05wyjb+9MdhylVvrksQ57r0t2oW/ofkfjoDjyqe+UOogt8s7D2Vh0BONk1ncPNivUqsmsnbgV
fceS8MYWQ5oE7G8M9lJCr9qaLemcgiEySP17cHadumagD69HuLwSF7tBOiSJnEJsLYQlOti4Ga06
Db1MkAC9yZ/sAPBbGr6JvZre4aY85kk5Nh5LKnwArBD/IWfPhFbZ7lAlocl+DSrZ+3U7qPvHuyum
R9VsloNaNASjgSxrWMnVZsTGPIc3m10ntobQ8lydZ3JwPXvcO+jnUOmJYssYjgSw8EAOYxN4hAJ9
4gzAhFJaa/oxG8xa8y/lSYek7aTTQtp8LoPzHizuqgAfOfjXairwGMZTJJaqhYe3SF8nsk2q5JVD
o1NQSNVF7W+Svm5/E/1CNZC166HaB9qMtg5gw3U+kkwo7YUVQu0nfOry/m3pXvOeV8z2if8s8LlS
BXeGAP4heho1CWTgF4zVwT+4ZgExRwLP7VizQYebnt4eWfr1QcMheUMMOE6l58U1+H8ppjiABYFn
HmWZ9pa7n3SAtL0U3x3Fmut91SGO2zz5OyrX3Jxi4DN3Jnjte5O4l30z9Au13Fn5V8sqLF/70z47
brxXold6rsak8YGUFNzLaucEeH+Z0yKVzX2iJByrmqfanFjnrxvN34tmpQ6p0IWjl+mMmrAvxN/Z
/g8tV7BitDE33cN9M4khevmk3extUSdvueVxAA5sqDjQm3G/Y7LpAuNsPpmSlMKDUfOe6rJuC1ni
1vk+WB5YPnXB9fYJP63Uzs+pchj5tjGCwpl8U1+s7iO7zzOpXhhkbv+FeONvmcbm8GDR+Rm4Ihvl
UgOl7ifeuJui5G495XBYS80EVI5wyqrl3C6L4KA8lzUQkio0MvlpKJ2Sm34YoTu/V6TalasO0N0m
ZuO/fz/MykBHCvQjLGHoETySliKmGP/Jk0Xjc5BK7ygekrRW/v6sBc/HLMK1EfSg2Mwe3anb2xra
w5Tku0N75KJXhrYc5EVHiSbWK2oN4d/4wQl/QW6LnlgCCh32MyQ/qZutmutOB2b2U2V25YOVYY43
dIi2bd/25ZHeyTlKlKG+dYcZ3vG+iOQ1oetBV99P3A/t6bs1rEqqdfnhB2Nee++YgIywYpXxqMdB
FadAtDDouVuowUO/qlzI/5Lo7TC8iCrYSLc2ft42xLZJwt+Ap9VCURQVo4fhwweHDFtDZTuTk67B
xvZMXRTUoOQA+5SwGPQL2QZniyGP5U2hRloDQ1eCST6O/rI8qCac72iAexAMuUXaiM1g8vE7GHD8
Rt3nXMQQLcU1Mua21mDK7OjU5wvG+Kq1sPmVvQ4puxuYUXHMzfni4dzaCD+VIPaME5aq6IR6ogpZ
NZXOSuCUbL42O+HxFIU1YWSxPMe00NBJglOm+fkDttaUEGxdbbaev5P0YF2kvExJTk2wAI/QhQU/
+HRniDPBwF+k5xP7RRot3svR266Z/rT8caOfYawklM78oOPh2/W5079oDfy6j8q0NatrGqtOLsGM
p+7BJLpxeWRls029xWJzjB2OxqROikV2e9hnTOuxbL3AGkXW2TcfMnLYMsjvoYsxiC22RXa0y2Ut
SVt8zCSrKb/e0masMR07eE2Pi94tKYKPF68WBE1MxY9lBWE+LSp2jaZXTh/6jGEIBtZQUKtz3hnv
V68DzEKx/uylCli8fclHeT+R6v4tC+bi8N2qg+RjUKmOshoKGVk6Qsih+hE3PdIxYbaJI8OErZDf
ONbjtPj+xkYYkpPFmKo8lT0hciDbXyiqWUMQ1DVicfdRLRhPSMwoK6nhhy89cU6R8Mb4Sng2m4Nv
nLUyURHGyRwtHXIJwPoW6GjyEd4WlL0n2B+bwuCqG+0USqg0zQgmBZo/u97Ml8zsErScVkgMIhzq
YPOD/p4pgp3ff97wbDtNSQkH8jJf/bcqRGnenxTFWGIox5/CmoFAKMSw8GlsNHTOBAE5er2DtODp
j3vJZziMBmP9uqdSTDNrFO437ufKdBMuSJ4omsnUOrAQRgtg+jQGGWlVM8ET4mYlK71k5tjYscuL
LkiVAIXxduH7lvkSsjlGp3MdJKUufR5di1OKHYS0AOPwZ02fhfTxSw3RwFHnV7IeniZPkgfBFNe7
S3GZXJPUwoNa3brl8vVDw7b2HMyVeKOPZsi5zb1x32hFFDn1MkQnFX3O+XM5iOY8+NNZzfgcSoWc
ZwcXDIuX+eZnxgn6JkEWM/+Pv14Dh/gbp1d8nBMX+HZ5H9b0TuB9Q+x00YbTpO3NdqRZcIzJqhA5
EXeVOcO9x8gV2yv7z1hCuUrP/E9tMwzixMJpY0JDf4VN/WhMAHwLejYJbF79fwEvoUwyB3EmOvVz
A7UmQo6Rz6MUTRMCiCdw5YY2+oExwZ51rJjc+FHTj+oqUHBmFKfhesXnROKDjpGykIMeHaJ6+eOt
v9A/CPVaJb5JdIEVgf81ZYgvidb34FfgH4PNcAg5JpXQuFFS0F24+/ZT2G4XIrA3TYPqm9lvtI5N
KhiZbM1jQRNI0XhXtyZbwwp8SCNd/FlJ0P7Pw6FTqj3qGwUeKq4qByiSnxpICvGvpjMOLjtrwSSX
XpZ4aQlFa0/cm1IdoEoYsXuKefMYwxUQJpuh2iutbkwSbLhgpTFvk9FTQC2u1s4plvuoqdYaBQpz
84O4WPRuTYHDvT9jyxNqXwwL5iFbzqjK9CaR66e7QRaVwfZW3DI2KOYHqIMcpXPsCzstv1oUqLk5
KV04rPMDXxMvujsIkBSp3TGnWe3s97ZpjD/tOX2FLbui+2NXOHgQHm1z0UCgEhv86W2dVcy1uybd
gy37q9Y5GmH7asSjAfeetKte0tx231P+yq3JocyeK+rQUiY5DcNJoBwfUKNlUvgeA15cuQ3OHOF9
pEAaky9vbV9Ie3RimHFBQ4R0vyqHHrQ64fz6/i20Qyh/EcOnA3WTjPcvqcbtErH9dNqvFyy+DICu
HOOOC57iUbCssL9tQEW0d9e0Nuo6QSQLXfJx53FI1wzkehV2lnG7oDdgJtsmARNcnFE5g8AR6i2x
sTNB/bgnBfFa3eJCqyVKcEvcOPpy6W74UdWWmlrrno8zmK+mamNqrDePIPkOLFe/3Kexx+nmqncn
ZKHLjPz48xgoP6dbagmLH9nEZ6hhIDeMeWHwRKf5M86EbOYJXqSDif/Hf0YRD/SuXem8f9MDiNz7
9IiqrJSLdN/u3v/wRvMzIkLpYisdNBpYMKW+gWFvx+21RVg1YzroCxZaYr0765aeLIyTSwh4yoQC
qP2+lIXfB+LbpfwZz7mezWJ9NE2m9GHxD4Nwma2Cua8wwA9MO1KYfk8bj/WO6tDG20D1eZuW2uL2
+fw+B8GBTt16NxJu74Am/VOcob6kdpJh18Yl+WuhVmR2HAwW4BDoibCykOw8XAnIVZGOBcnUtJPj
2GJgYRdLh3F5ykvgdlXls7jHVSwiu6cdy65S1PSaL/f3sahBPCkPQLCe2Z0VwnGMyxeWwXY886eb
9RiqsB2eNdsChgD9fVzpTvxlvkCjAmrq8aBK6RUNCl8n4xpH6hsDu7uJdrj31oXe0PiNWc7EGUpF
XQ23qihC31NkduytPQ3YvjkYvvRxiB6xniOxpAH6iD6+UMRSDwQ4N01TBlQ0PyD7NsxVrkB+FdnF
mdQBfLmgO7faW6XtgDQ8uaJeB535XTjrIhgcGDFhghxv49GMBzWYm7hhquN17ANAkMcIiQiEQDST
Xs09xQoeU4i4CqBA0tkn5rrZQAtcxMXMJuZCIW4Qvw468cXMBTSI8LdIjcpdmZEyL6dj+m7uSpgg
5/M0LCxQ8CM6ueUZQpkAqNSaBJZtgeJ+3Fpkd7b+xikAVVyEAE7kNzyI4N212iK+R4vKTy2YZ0Sz
uA3ugSKENcVqthvXWDvxnccUcxrtHbPwWAvQLFlkAXFrK/mXu2/YhqSYY7tPJypZI7qUvzBWZRNs
VbFgmT23tFvRsPQVnkfPA0sz+VVFVURAE/Ni9BcMMgq2eVrtYNgKb10vaPznzo5yMKrB2mQJkZZf
CHzECSuYTSsbCbYrdeFDRlleNKxcw5FQZ2AZ8C1RbdHbXEyJaLUtDtW6e8c3gOvd59EDn+z3PYva
AhDE88mHMCcDfShKRH8P7zdAPbf7KAygVOJAmaiz/i42OPGQOFegUkFqYEwuTZSn59GcM7jy5SRl
iaF/dGlvmOJuA/Nic28HqS9YNPvOzOEuLk590Z2CV5R38FE9M+10Uz4/hWcBcMAI4EqwhIUvMZln
aeJ5UQ2kgqB0HGcit9B2ZTUsBpy7CME4ItVwNz7U+3XiibkMN18Sx2b87Cnr95WL6FkkJsUgw/3J
bVhcx3GZKVk314Gfv92T+ptEmInHnRlocUP1V2Lzil9qM0hSpIet+8LqA5wek8yHDSz5T7JACb9G
+SfPLUWODvdvIS/AzhRmsVxXi5dAL7JeRxErr5euA1zEIwKw2xXX8N53BUGH1noEsUuB+ADfywjD
qcAHw2qwRvMsVudKtNVf2LeFMLkzBnSaBsr+yLiI7ORFukaC6JeWeRkx46VW6lPISyhjkhOPQuD3
TxxsgSNIhC5NMm4gxnC3ImXtVwfXdB/Vh8doYzMNlptKPS1rJHZZfv9p4nHJ8mJfWX6B4NLwFihy
rKs650QsTsG4GLqzBhCxiJCnWum/RVOu4fU/tk+42g2CgaG5BJYFL2HzkG1yRxAbziBjIAXz27IX
v6EWTwzUh1R7I3ecaZUE2sUhkFk89vlDz+7YJMGhPAMFwzNb9n5FuG4p6o0UBeP3EpY7vrnb7cWp
2hAdWuWpVrBHCMDaGm0C3eSi5yoKafqrm4GAjd4deTmDhWtvQMcckqSssOJY7uqbvEG6fhZDFf7l
FGhN2G42wj+EDZq8M3vTibdCy490KMWpjjZp5D8wLtqe7VURB+2mL2o70fiLK92BUC66/3OSjAaP
VXUcabX5NTtRyJBcEToqPBzfzp6F4yKbsHKlf213r3v32xkx2DhZfdA4GX0U4fWakAuU42zLzBTo
Ede5D0/GofWsugTM+wjYAxB11Up/arslVu7mlUrSrioFOkscaOSyS/lXR6E3WIubkwpnk+IyTpu9
jNmPxJR1OxmBwNm3wIVKvSrm5PmzuEZqCfnUT1amITeco578itC/IrPRyZqBihegGUVICkDLkhzG
mz2UPb7q+fwC9w0lR80ua3CuKK/FTspctpr7J8Mks6awTSW4txf6u6QSE+wy7mi9ciR0IQAFMQi+
BAYo5n3bCxDel7xeTPJgL7yNHVI/FcEUrOwByx0I1YLkaIkdn7ogqK07FVVCMeuiT0L5p8Xf3URB
1310sE30RY+lzKS8ZJJGT3k7XJJ+K1oTnE0L6TUipiHBfkdJeaF+RlArH3xLVVbmGv/lkAbNXWhC
xxV9JAjoCyXmCqKjk2p2pIO9W21c+R0ydrJe9auvTA15e3PAhi2uVHq3U8Ng0IVURoDvC4G9KEYk
/p/kmzmhHW/F0St5TUzLeva+bFqkH1ETcCTvVGQZJckLQwpD9LpLSAmmgQ4eyreNYHCVfQHf3IVS
tgWqyBkGNQRN/Imbh38BBFHiG1DNEfXv9I2WuT00or+n+5NR61Sv3qX8TVl+r5pbc5z7AxjsTphx
spsQ1/CMKvarN3zwHegZwnQZEmMRsWFp2mRdZOiM5wms4TmicyHri8Wuq4yB9qBUYAuveI9ncamo
7YOaQgeJcdys2F4vqr7PPJGYTV0eAJHSdCkDw7FtChlfB6bQ/2VRXpzYpxGDQ5b2UDfdvsMqCkrT
rB5pTsMrN1GCiBcVxMUBlNS7K9R5CNmnfdeG5zxUyrssh2ItaySsSquTGpeKcY6/8/oh+QihluX1
6VKlm3PnP49V6PY6H7HFmFr+YlCBqyo/fMI4aVvOhESycPckzyj6I/lJny5agu4M3oT06u+LCwr4
GBuz4cQY2i1pA4/cIinmQvFImWimp/0ZAql/LpNmmuMLfWBK/P4B+pQ5qQHYJZ/b2zHyN2kxSCEy
WFc78O7FP55VcoWjKwwuQW5jVEgfqAGd/YLeIe9t10WZpneZP6FupaBXNf/AdrTUJRet5mCJM95m
20cqicGXza0M/Q3P/8caQ7VOsT4VMme1rAfxJz9B6VuNUf45aUt8NiRT0W/QSQD65iqN6J+eQMww
lYnM7JwL7EnVnMiDhMUEFkrzJMLygzpZKf44WE9auV8Y1Kn6eInSLTG7+C3PTOWjqmDL5bw5XEyg
AcByA11j+vGjGk28pydnsVPbXXwWRfODn1dCfej9QOVar9J5YcufDjUD/rGurr3rgSu/nz71gOpv
iSfQfar1iuylxNK/8JH/VXNtvOCWVmDTMi0+VWwqOgeRbcGgUicTkjy8WFvI4XbMfTFadESKqbZ/
nFGVDuXaBUnuxazRmhFdKJh04ZuZRavMd7KynapkePZBUC9WutxUkti+Wq/9NCulB5pbXus23mhW
pa0yVAqu0lhIa1cU9TSEyLu/LqxGaXrw4vsB6xoUa+LIQTBsN6ujyVesY0Qaw5+dxQI2meU4tSic
U34hOAIXGWcfmTrL/J0Qix3prakiV9R9udcMDySVr+FxCWzAmdaQlN0AT2A6ZTvvgOA2GOyF9GXk
sozxYR9r1u+wMcnM69s7C4uWcaRLPYhfhESXL3W/HKEUcx0OGjZcLtAfnGjPY6PfxVJ26ftpy67b
OxrNHbv1DbVtlsVytU6OR5XVBvqdJxhLJWpF2Qi5u0j5LmyNpEV1scN8SY+J/xggk51P9stTvUAO
oEVk0hY83TCIhtDrav0eWrYWU5yR2ipYqlmQkPMG543sqxrTrj/fAkJ4EranEqJQ4gOFC38lmgwX
2bV1VKuX+c6dEupxa4/O9J2I3el68Qh3Efwx2TeCURjcRcEk1QR9f8ZctHspTEg2UxjQhNDStSg7
zoCZh7N9/p0Yu22yRbM+GY1+l2f0vObQcujbCewIHfKjvo4t12zT1YxWjAX5KL+/DdoXaCJgw9YT
82X5CGG6wi/nV8U4PhIapLA9RduDuNz3SF1DW+5L67HEHOuBj1BhAfavL1URPlz6NPpyIwFO/n6W
kO8JvdntjPoTt/FPfrWvmxj41PJCZzgk0mNQY6cpTxLomVCcKFHiZlUX+BsLpzvJm0X9gGOdzgRl
d/ZlkKBwOcP0t+i9fLGi0fWl5HYnrZEtFLtYmbsIiEGWdeWOK2PwB6nUYcyACg25oxUI9l1nHerA
Us8Doz0K1Qxojhz0+vYbozczO9RECEt3uM8tIAjJDIy5CeHSSAc9ORruvVStcSm7VEkFEMH2BmHO
cna1Cno/SXQ+4cm8F8zmUx9wNs805/w2oOE4UuUprSFsTyEnTrB480cYqzys9DFRvJJemCEYYIzx
4T6rxeyHq2xlKWeVNeZT3uIIF6k72g2/3cxjMocidgLhHt/Kzvan6eQRkKni/QpIIEH75TdGDMc4
3F3nKPXzb4hz9vC1XUsxRSkzBiBVJt7jreSpESLmbd9KtwHH/M+8n22hrI1yQBfFnHMFldrCyGuc
8ezRCCDepBzdjXIz47OsBCuXYAv48UtWt2do7NSdeDLc1I57PTEMm/cYHAF3/klEOnxQo9Gy72nB
GrP5+LF3TBkXsq44bjZMO4fm6eG2km9xiSOYxjJuJVMSblVjA24UGjlosXNq4frgpEs1cAD/2R8B
oNQOixTYtAn1qV5dt5dGXsAqQDxJRqXPcENnRVCWzmmpodIx8SzzheXAyJw6vSCJI3cwuKIprZcO
jcNTTKKkE/QcuB/b8kPBPGEahb3J4f9/GID9PMjPvHndcMhY/6ouC4UanYLeMw2bDqIKCyjt5y7P
TNX9V5U5bmEOVDzrbTI57hG482xPs3iw57eZQKqzSFpvQ/yfdha7cye56JtJz1bafVy2RLTqzrF2
/Ibjp5QAhZHABg3UzYFRcM5qDMgkAhMQzCiBdgRw4Ey3WkH1drcYw1jt4fKBZvkrCRXRLs9oQf+R
2bQzK+7HCU3cUSBodRbte241IaNayPrSsedQr5qOem1JtfM+XXQ+yaao46kW8MN1M9RYn5I9Td0w
2rIGzgxEsZwDp7uMWZ3yUBiwj3uhiEGmyXhRXg06qtCQFHWo1cKmY/6GzGJ7M7X285Tl4Ml39ZAz
W5LNr7W4B0R+xNmo9KjNZU3mZRuLL4O300OhvN1Q7RhtdzUrb8Df3XCYuKdUk3+s8Xp2lVZM/hFC
+4PGD8UUNcpLabZLvBS0y8AGKWUGqFemTs0ZcT0za18b3UnbaK2ye8XApl2PTaWNXJoJ990vJHPP
VQwCqCXsGqWfRthJQdTDKEDjD85ftj5UYarNOPgtf7Ik8oyxAnL4aW1DM4U1KrAhyWI/WeyQ5L/W
8Q0OPB79rMuRasi+jJb36c2cE+9iRq9hkiahtGQv4w+D2xaq7CoJrUgvJg2XwBKmy4L4I0ORMHkA
LjxQuC+mpMzTXjZUB053C0CrUxPmziRdRO69xFVHBjdFLKYHZyIim1u2z2XEASLsnmrU4QoVASPj
In1C9GF9t6eZmL7eF8ObP+zjryw3qguTM2FxsaaJ53sOuTtIMF6csZT+BauqtDCRxGWFn6hRBKZ/
Kj7RbUmjYozaz89T0uEZXqs2KTT6d63+hZiV/NCvrXKBGQ1Tt34hMQVI7D3cAWoAqT+bI/ZDJG/p
dkmP4y+MaP0xOXigb4THYBuOOqZ9AniOeb7H5AJeOYUvTkRxYEM42eEk2c5HyVTi9KNjVvQv32eS
MkwtbeJR/Td/6RWFs8VTJ26a3FvLtPlGAttLSxJZEMnYPgjDQ8oGaZdIQG66QpLKkSUqHlVUVLZH
U7Xi5TVTOffHjEHjdpl2OBCk/S+bhlEJDHSR8ka9pUPchNQ+vuyLFAIS4Y/q9tGlb9z7sh7KvkLR
317nPzOrJcNQ491ZkGZvcODXA2CJFmpkBdojv59E+m6GgH18DutCshYuS60VkwfecHhKjPE+Oekt
AuhnSJM+yi/G6Cn4LH+Gnu6+oQHxEmdL4iExJcvDpL/8KTNJm3HqEUrbf+vcWzO2j2UtgIo8dEPJ
Uvrog2kOp/Ve/ypBC+wxHWBfE5HytPqaFG06uGh3dJYSB4BvSyz5I7IfGW99YiADpHUoGAMc+jir
Bdqh71mOCyEcVISgqDDekpeddEHtdNWhgOYnLImERI0Kqx4+Hl0CqY7H/Yrcc+KcnMYgLasx93Ko
g7IzcOmOIP88xUjvBVrg5LAkRXoGyLQ36upMQkflLDFJd0+wDId9FvC+NFGP15sk6XMvdcykYhNW
+50CiW93/Ri+XNoFuZsAClG/nqL0zuZKDol9g1Eb3YLuxe8bjKCgOYyz+nu5i/nqZllnPQIt92qx
B1IGLNLa9423NAXG8FwOZ40iSQHh8msh7waJD4P/EZ/nDsvBC2iEXRCdgmxzwiwDY60dybdh1ExY
kmcSSNTOu4+jpB1rleCTggoiIXxGfP4CQu7VEP3YUGkNGogMgqeJpKF/Kkqvz7v87qri0bN0tmmA
sAgEwdsgDXUEG4lk/WqJqe+2vQZ090W1InAzgKken1AFxVB95BsWjMuhWv7mHdKyzVkwkvMVWv32
JFucnLFIrRGyxUDUJ/bIrkAwGYg3xtOurfl85csXcihjSIMjauV1UK776U3vytN4XMvIMrGG9Hes
ToauGrm7KD5B7VS5mOFPMv8CX4y1IcFlkaFKYgbFdfTLKQzBwNEdAvvqtW2mfZeWSAhBP5NoXIIG
2fRxrIwKBwP649Xk/DSqz82C2Jr1mQHtqys0Q5m+axM1Kh4H6yxpfEYmFQCnRm1biDcUnLpN6maV
M+o8RCkKE+9zRrJ9skokQ1ZB0qPHG+m0l4uxX7kpjiw+FQkxw29LKagEoW1HBd5shqt0h+ClGlwU
Wu8bsPu9Cjdd07TWsLvD99ojY9I52+psmYV3/r7A9gaP7mSWgktQnKcxJnoF9sCDhwcu73Q57a/U
ugOtxMzfsp/DWOasUzc9eODZ0IuYqUajS8nFgxHa+39boQxu5MI6q6i/0EPvmu+Sr1MePX8COnnd
zRV3EicmH7HVQeze15Dj7LyIzTInI6EJye536i13LlCrtFpLSiHhOjpYRe+jCbfVFX4lSxuqS7QV
7HZvuR19rcHwOthargcRTftihmEay58BXwgrUXscIZuqLx/LZRHEIUubVRAF1D0kWlGKLUUCmUSb
CErHd+AOnf7m5914wjA3xXcAONFlmP7tVCou7Yr42MrMEFaoWtEl05mbVQNjw4FqN95UD0sCGx97
YMp2QtR6DvrpUtAUAFNdJl1MUEoQWDTD4E/DNUwWyJLlqRlzjO5mj36vZzc5pA5sUKgyoRZAkOL0
wPpwajp1gJeOuy8R1Q8GDzlz6GJuvN5XsunLByoVyjDBtKkMN2o3OcZepX6kxCl/ETpK/4VXruUF
Ze4HiqS//9+9SWxT/T/WC+mPtSrD10I6EaQavX0ZdOVRYWcS6VZnvn1xsCiytC3R3vFp29hqoG+B
TPLum0u+qXf0yrY//ZCHJfMavFixWeq4nI7GaLukEjQp84nqe55QypX98qYG23yFIZ+WXj5OaseH
4/Fx8NArbHHmcNRUqTv3Y5fDoIXQvEYQ1wim5j19hSPI2JXqdhJOiFfCaHJFOkW0+IJ6AQyR2TIq
6xE32+qdZ7sn2N5rwgsU41N2GobHnrfiwr3m9zeQlfdjO2OPK4bViI435zfqY3uIX5FODsA0ZLbv
1IzboK4isp/SgQiHu5Z6VtqcFUKjZLp/JFvZFuoZ6CApa6Q8AbAQjT0IWcKAGdsKcTloRRFwVrvS
EE9zWPR9UX1ybQlEjYE62pzmzmrgJRet2SXt3Y/Jrf+vAMxavpm/y7BCmXlMN64IkINIpq8jAhbT
k9qI0wupU/PoGNAMCRkn5dGeRBf3TxzAGrMfQwzIbvueR1x83Hjksr55zIB6bsdANkXb0ntv81kY
x/pcEfZ66dG6TFRDQdE84ePCmaV2bnOeiu6+OQgRGV9RdnL1AanWzAvzltdjdFRijGCLckxSMAr0
ppLatLZRAsefs0uftwZUvYfdl+8V8eaq9FxGXgdl/iF84zQxKAgbP87SHJ1NIvCUT19svkV6kKll
eUj6+eaVnbOVsYzidIn5/jKkmr2WPfLFYLGxgWGzeZa9aQovkMltgqmeAo6ZHFmJy1v/b8U0KkFC
7JIg5bPpThrd6IjrWe43vt58SIeysV73b66Juh9WKb3/aMhp03TDjqqeFPYi3iagZo3aySoOjEdY
Vz8n0yEuX6qFTVAtYNBULJh/kFlnDBqTp2stsjXxBCXVJpmsKZ893EkBkG6v7NWobMzyL4HPUeGm
dQPVHaoKvmGxr2FVtaFFaq8EZuXvafmw0TUc4fnEqmbwmRDA6rl3lq0VMSYJDLFgxDMpsM24F1Kp
DEtEXWBkTyvnAZM1WlsKkOLy598d3KFj+vcL2pqWusvAuHCl1LbxfK3+7dOqe3vkaiAkG6GonAoV
IQD//4YSriFXAAC0m+XzN+351DmoxFLDOjAspaBFlIkSm6BYmqVtLS3fPSlDDCqsWptz1wrGu8Y0
cH7OW6j9DWM8Js7WSZX6g9ZTYBAHoDBMP12qb3fxhksFIuCo9QVUvZ9AYX9tNHU+SupSzFwJyiLC
ENy+gr2DB5xvCGfdjdWKcYHu432/QbKmvqKrZe9hbO3rg2dM1zZUF6E49AHApTWs0NerPo6EDZ+Y
2sGIdbAirWxf2wV7lZdO9FeuOJ2/7pHORb8dxkTIHpsAuLoLEh5Kb3MqFMxZxvvjkkYmjodzmHri
NLASImhyTMYu3Ac0Pao3D3km9T6eBZD5cyhFGw0mr0O+uCWA6eO6u7eZjNULyW5MnzEeCK9eJG3k
0meXxM//8GjCU3njAw5CIakx0OLcyKcPnZEhZk8aaVly/QnIVlmkSYRxoim3PKszr9bWLDM12RML
2YiH3jWbxcMT0H3zzwEIT9QdapspIffLEJa7MbZE4Gb24rqB3NzCqP9dgsyNuoV+0CGPcRP5EL3A
VnPP4SlzNcftRet7dNVKoW94UQvHuA8z2i5aIOyKWLGtsfeEgHhw8bRqbrPc7HmVjne3m7gBe6ak
6Dd1uLncR3p9VtXKbO6QSdve28Lfbfg/5QlIzQaDFX7O6w767UYQrHKsx6V7+sz++lhz3EfF0t8O
ZNAamDw/SJbXfhkpmrJa8dxp2zFaIuFZ4yiZv9rG0YDDJoGB0IBvzXfbDfEfajpffsbOB1cLivMe
/MQPYVAoqs2v9l+m70lbSUAkNse9LoQ7/JyOMpVpCuOhNnQfARkyUnv9h8iFhAPITySl91hH8llZ
ZI98qVqW5raak5mhQP6mp7kJ06mllqRpLhklW3O15cX5W6cqaJN5aGr4l3qSRaYeNaNBAqeKVf+G
2Soptib3xzcMe/GP3xudlwlLZD5nsMLtcEerq+Lialx9NrZflpyyhfJDw5sdSwOhoARohG04IFdj
QHpYY2fmC4Dd49YnTUg/HiBLjvhRhUe2MfsBrXEuw7FDQIZE3hnheF4JXrdQgJ1A3xuGjqD5iz8Y
8kx8QoEzP3d9GhLM3CgdWu6X045DOynqPjetelH/QmUdeTlnmJiOcjG4PZ8mrmQUELvqDt47VNb9
v05OuuxS+Fin11gkr5HnJkK9zHribyIzYDjyL0K206E7+i4n5aefGwT24I9lkasw4oqa6pJ8abuK
yoslnjYlgTt1dmQMAsHRBiA0MnAjt0OOUhUd8jZe7HTZBuESpIhLC+1fRXvax4t5KhCjBWPgr0bK
fsrG2YUPdTtz6trPZEkSILxMXEe4VqH7ZH45fxKHCIairbOxvqTo2P7FQbLaPeHBNAtgj6he3b8b
TBWle427KQC3Jfkrs23I7jARWYOJ8dwVg7SnlE+o6mX7SnIocTWJjZDTvNdPvcfUygv7eGmcZG7a
fBQWTvmZg4uxbGbPPxA5JHQOa7iASn+QqsL8Ad/CwbGE9LMrDce0jNVSDL0SiyEVTxq6jujMLkAM
Zf5ySrnWg6FDxNBPnrXirs+ogxbJBOA5WLykIzdQGGgPdPh8BbQTfE99uZsH+cGOIw93NvTn6l3e
xqUUry+8BTfu4oAh2xTiomHCEcA+MkCO/zIND9NYnyDGawgpHoLrtT2RNduVxyI/d05U1GwEgvf+
O7rfEOU/vLtMt22AAMfZR7VOZJIvP8IJYL2wSg0jkbRLlmPkU7Vrq73PlWbUr6qb8H1G1oxISL7O
HlQvjQOrSCC4wJSDKdC8Yz0xPhgh9AQXqazmFcE6M0FWM97DFkC//HvnebydGFM7w0x23DV0QZTv
i4WxYVEhkZpNBjX6YVgGX2q0V4j+8szAV6rLW5SZSzA7TtJaYB/pfz3GJIvJYBCeG/Y28UFsnhko
4a7aV9VqcFx0ufNyuio2R/icJ1QKJVer1fuofcAomV17Ebu51ESPEGKnJIvSqDXgEztkYrKPWWOS
Wkoz6fiGMW5chvaPKvE3UH8kEgHbaElLG4vFqGgQyCnM6BSVPdLnIUb6jIJH8+yqIZtLt5ag6fK3
hdnxY6rqUSgFOEhBjxGCQWqS7XlkXAJwhdoahbadEY/Xn1fbWP4uKkbpHup3pMDTvagUFR+3fyw7
UL9DAADpRACQTiGmRA5hjpqh6Do5GhP8pWuxCvcjSLT1ce8SDholf7vYZrm1dCYtI0/0j1og4WIZ
EyfMIrX1kraa4xJGR0Vh+X8BNNQcUOiejEgviaGVmG64RW8nI3tozjRoBtiULsIkbv0+gI9VLwWc
rK7UslNR76yHWEEps+kiOHdYCxB+wTIUZWYX8rcdqfTSwS5PY8oiERlxS67/NDcAxHTuWMw2Ga0u
R2NNxX93gPoa3XkFuTaM8vL+C/wxD0r0MTr6Rh46KdnVsD+e9JXNOXWrdmyhdVCFK9Hyk8v+46oJ
IB+lHaIaZvV36GlL5ISN0YWHny6wF6Ex3+15+DzT9ONy6clmFDF8abbLGwyCoTmzU2ogddVYlsFA
4+iLZZ45o3NqsPDhbkMOAc2cC/k1AeO/ydl8IgbP/q6TLgqbSyvD9PvK8Am6fXPqmAme2ueP19Pw
TQ2oV1MyvO0M4I5Uc/79xEwZcQLVSM4DRSsWssZ1MahbDJBZpkeLmgnelNV0sA81VHCUnOuSmGRP
u8W4zwnbSbtYxe3ED5voQmK1s344hEtJ1ugF9EAo4uE2o5SFQD7OEWpka6MHZy5OjmS/8iWnCuzP
0jcI/5gLZZaW9UCfmnY2TSp2gl6hdorkYI0wzf6Yia8qSTiQk0zcp1cOfSxNjXjIHDTUVQdTRRiS
SVs28Vpbf35uY9+WGx0AOmTkNRhbaLz9HThFyTkxTJzwkz/HjNWgkBXaHuF+qhCRGIytUBeorgPj
CguCkZPPT1EWMHcNe1A6Fv5kMwKsJa9KACiZnSd7KAnVNdJY3KvUEGyJFQl6m/KXWmokeyBIPhWK
lxWGn+iRNriyUecGMmLbx0rmxgz30Ad0JyLgXufk056QJJ4zQr5IBJJobAGh5Pr+fHfGITwzTuji
oniwCLMKKaIiRzcukyt3CcfHwnZqdt8/EShZEkcuT1RMeNlV+7vJMDFQEiATLoFUqNfrvHNwTdSY
mDndnJPBx7kcs8i6YnYfFJ5MKeIh3l27b8nxkzq4uZt7/G39R4H6GsmN/yMvkGdU0GM62d0A1vUh
OkLU53VOJKMjvrM4F+YOhza1nnT2BAsLnALrZE/nNIoeCDvyR9uN6uAtlHLtrYLLTJDCjJdYul0q
Owv0ap0DGq2/52ZnxMlS6O2lqFhMD2roMR6IKD+JauP2D3kaKd8oZSPPwIuGHxzfE8I3gsSGntc9
y4Y2tw0qGbhbKNM/dbxcVtNQWlGS5kzcqNOZ8BDdG3lPGuHsobXotUS8K9nHh5kVDsU9KDEr5ryr
RYFzmPKZj3xe+6FAoDyYJQPS6dUSw6vkVb3Cnl5Tau1MJTGub42WxYf7XUyJwr26jmWBl7dJ/x9E
4udOnBgCOF8J8Vbbnisdz8j3TPOe8FIIVK2lgOanCRslr5ccWHEw3LJ0y3p/P9eEB4xPyyXiNMSB
vaG9A1dPaD6M5c70KDWjoVDm82aIriDxQfEbfrEaUnCX+IvmBNVJnFitX9AjhI8Z6eYVEkxH7X1v
jLac0ZxDK0OF2SDkIXRn/bVuvnmb/BYzMe8O8Z4dHTSipdJmgrK+hjYFyXZvqYuw6wLYVA4FVy9D
Uiha0dQm4oJJrk0qZkAaF86l0fx9fxGkWGwYPJSiX7ThAEtyPgJ6cT6iVwedtoqCZc3mAzk7B0DY
p4Bskj2S+zVOh5pFXj92wjVKUuY90pbokAxEtJorS4tHME7UzHZKSXR/2OonVIH837dXXMb/C4R+
MQdjcTPwWRniz3+X8oOx5bUl66ClB9OqABsEyhBy4wfwCgW89j1AHF1ubjmz8Kxz4n852E6qfleQ
VpLABVpzKOtFZ8ft6PIuUpqXWdoP75vErZefvKc49gokMUrfrWrXs6EMMx5nYJMvKe+ujuGnyYbh
uw+8OmKgrZbCG10W1jFrxnDEWKwbP4ZP/cHqB4zDKAvy4PibDRfyHNTZnuiL+v8nUFRsZJ765MrP
dpAmtmlxyNMk1suBklZ7kiNWKNs7V3APH8pDmrGwAibEog7cxZQ/I2qpKDLlyPCBK1YLL2eVu/31
9gaiBHRXn6rA1B23i0iLleWfzlNF6OlhfKNFk7xtfZoz//ymJp8022I6EuS3yWTO0FBdtU2BZctk
v5GTlXvX28WW1VTQi4QmN81ywO8DLC6WQ6HF1WQF6KSRM7Ps3ica0mLmtFUQtKOuxgSlsOANlG94
p8vgc1P2TmCYs9NVscNTcsY1MxpD1kanW/nAtH9zPiM1zEbc+ul/HVkABalhmFbV/4EWk2SHvUwc
jjsnZQ2wOozLANJsLOADPcBawoJAGf4uoBfl451TNm7jPG4KUI0X2+XhJpbqY9wTlQ8vxTLMkgsz
NlrZngJDc5BSTPSta8E4zsnOR2rdvj+cijtMkLeXsPx3ZCIY1DYjvSza0O+Ind2XA1ZQF2LvNkQV
dUWk/5d2Y2OiICY3Eq9Wqww6gxXxTNTA9lZpHixtYq9CRq7JY5mM6mXCE+AZO7ePuZPLrOetqxeo
+CBAIqTns9EcxXIj4MCj8MGZeO8xezcPXiQgfSw4z7TJi3eT0Oa6qLsa6oY3vUr5cbfjtrOiBeQS
mKQR9lIT06zLsSEH6z+qWqwi9kQI8A0fyZkR5tomBpsCbLOb95D1AKVIWf/3MwENaAvuSeAvUmUZ
i2xgamG8VAsDBPiIOclayUJoEBwso+xefzuYSWEFcP7WSpY/irMD4c6XFGtaWvZ6bKXdyocqSSGz
lG9j4MxBuGkobB1TxEHXcu4Kl/QqTZ4UaIAD3Pq8HgGUq13TrYRTTj83BMfnfYLtnyhRgzTcR51g
Ds6W8L7TVd0iIJtokQqH/A1gYGv+j65neG8oe1RRwoDt/hFLf30v+L4HHiyuxgkJT8bpZwM1n/PQ
A+xa85+nShBL7JOzeD4eJ62IEwHu3P7U/iZ1fhoAELR+ybf05X7UU9RQsCsqydfSdD1q+6o9hZR+
BiPipAJ9BD5s+94ImEOjJrZpFF0PlhyLQHfJxO3RyNgec64QE2M9wdhK6l4y+Es+8tJjh6MjMNeb
NDJwSkWr9tLobwoucp8D6vYc4qUswoWO/W+VelFIdq322DdkL7LC87MzAXiAORygwu3mTjwLjtjH
TR82FrPZZWVmY7C+oaS5R5DOK2YQa5I+l2C10IbyskSe97/PQ0GeoEvEWNHMH5Nf4Bb56Ea0+pFH
UjbOp6HSbrpR0/yaZZEiLE81so8iN/ep/6+3nunT92GnVRB1e7qrjENqYx0E7N1wSjCLp73Lx53K
P0D1lBMK257FMP3S+iM3zhspxW52POx2PuNQ0EGyS79XotsIFeW45ehKFrhRZ1SyCrjeQaNfGPCy
WXvIrr3lTjnPx9kgSoedD4GbJto4A/GU10ZtonN3407c06J/cPVohtW6p05kj6yjl/wN8vieMwmk
zhC//vuqb6cUcN+2LAxEX1ZFxXJoi6i8MfR780foN1cxR3ELwStDtGbtmmVNUgHvmheMLvzrNjLJ
m6tZP/3AtzbS8E7tDx073+pTyozD3VrTSwlmBrJyQsUzjQG3Ts0s45WHCD8PCQIza8HTI7nG9/GC
F2fLwxTnmpRL0EpJ6wYiDbXzAH07r+Qjl22zvQQ5/fcquFZySpR6bzYwaLMyKdbIEsXDSu7wphJ/
yudSJ7lVAFp1w5XLrkpycbUCJIqh8P8s2kj8pl/0pfTBvuw9mAJZM0fYFNHiiLz+P/Oo/yFh8wwU
PKrw7M97f5Bgct6YEL+H1iMPHcixJ3+cjClNsDpj7CgiNTpvJ6kFgRsHlKrKXcg3yxwKtYFiTcix
dMTLEHs+DaQlWKp1ept6wMYAhv9KndV2tlJHxGgyld11LY8HrEJ7soJooL2CGPsXczQBLCTQQT2a
kk9Ou4qMSQx0oHP3riXIihjefan5y9bm0V/Sl9qDmX154o5Jfw1LI79jtMSONviJUH9px3uhASz1
mcURehOvOFhvgYi6KAmCLf2BtkomRnvxS2EmC1mH1mOAi4XrquhqObcPUj1GjzJLvSJSV6zVJcnD
ybrorymz6XInFoavC6S4+GkCDMZpuhjyhi42B70AruZkfsmdWnHrH36RXnNRWh53YPF77KGzYWsO
LoPJeEu++iDxEWTNSGdBmFr7pjbAKgKc3k+Gw/2F4++drnD4ORq/rnLWtLzArXOuNG1VddXOcRnb
ncXIM/r2hWrACQKnw8HjMM7HuH3lrfh18VLLfmQSbtAyqg6tsgWvoZHNSMIoGD9+usk+nrURkan/
Zt09h2GTK0hJYf/Bzzo+gQXYB2MPpsUUjSioCWWvzgsaoj2jMGk6QZwivtVSPTC0Wl00DOCau3rP
KNAxAzcDkoZxoDeR50nZJf1s5+usjrpTjxxCLOepxXvNg7fwBTNKXCd6DwfPsWmKQyLp5DQH8tkE
h0RRiarHORevL7xngoSAIt87Ta66+IH5CCCHwUg0eJ+r8Fv3GVEU7OVOC+rimIvARstKz/MKv05T
7aZUqaHFx8XltUSkep7R2Lv6FxIoLoAk+N7kxraU3pwJv6VFTI5jlVy/Q/inKmZCF7m9zJ8Wd5gu
tGWNc0WqvrSQaKfDXpjyu1DMBc2xHj7T3B73RwNEjQxIRWWrIlxhiW34ZhF5KPUEPUiEiWF01COb
SHA1K7noGHRIRzshGWa0rQHvuZvuSmHM71nROzzoNhK0gALsur1aIQUBfE6bQ+V+dd37kX30VOb+
ycvvpa3NOxOFgvWyF/gBeEgVB8XyaESZmdEMy2JVIPqIn6qwIQ0xmxZqE1IhtWeOqWbXdNKSNblO
rtLw+//tmye5hwqXj9FUIEr3R1fqf1k7hcfeUBRdbeLp0IbaiAwEGLZkhZpqsvIWGVXMWAfjKrZu
rJIXSle16Cu6hRUeerw/BWQ0v3Tc/WmaWx2dhkcAIHIP52tBKEIYPG5ONY9BoZDd+eOrW180pil6
Ced+UD5ljIJJCLmuk+P7N3iLK90LyiD6KJJBzW3h4SU1Qr/06LLHE2AYPfa+uzZBwBQsc801hUMw
XWubB/IxMKAfZy28EuKDfOGByhpT5PZMCrhVbWYHdel/f7i+e/hkCXsOwRExpdhkggoahYXYGUc4
KEHq9tXhjlUs1rQ30pCnyEjToWMvEIT8WD0FE77mgT6adckvETxqAYJVge7/JzrEJv9y/bWe/1HY
ZqPGbdGCB5acvMz8ESglq9c2gxPHoMklKd4Zqqavh19JbIZ/AuraIe44aM5zuyQ+wDB1b8d7wdMG
iBXWvs7o7HqWQ/CmpeGpI2emYPAojHvam6ne2sjUAS0pKrt8U2tUK+5XaHVq49J9XDeH+J+0S0/W
3HARx2bw6fKi17ZJPAFY2eyU7PFIrcfHc97lC76a4F0cK2YwFJZgQTnBrstex2ytfqnK8q2HmsZr
zhW8rpNr5D/fg80zmCUtPVpPp9ikCR2IDp+wXluWFiSqvKHqIjNiP6OUp8GxcH4VW4O3+66bTXgP
mjt/keUho4AAlXRSjyiszMvfoNbpyDuGf20DfTL3to3vfdT/pES2P5grgWe+R1jcse4K7vJEpQuC
zs5LqWqbabe/XEAnoysZ4Hiwm6p99MC/XaaKdsrK1MDt+JBK4bNEdYOws2IV0CqDcqkuJbG1CQc4
8Q1fXKnI4d3FuDkFPmmqzUx2qkQuj34d6bXlasf8p56rjzt5rfK92vpeWFPnvaBRjq40pJnguuGH
HDbMAFiFGytk/cGgJOYyXUSE6rStD66pa+q/i/F4X8iq4uyxUeSXN+dQJNCEl3P/CQvAyK+M7KlY
mYbZ7OTVvMC28FPzd786gwvaLA9ssca7Ay8AuvCn8+CW9Rz6p2bnZ9NWAtK+wpy7yf1zWOcBSUQ7
YEKHpHiP4UrwA0eu0s0l2oP7HvlkVI+dW20dEbT35bZ/YE8XhD9wrkwL+uWebqc2zG9WTLl0hIHK
wnziQFhBnTsiGjwyo/9IWbisVs4FfJrga6AKfpEGPsa/7eoeUFt5g60tQcQbsmCyVQB7/XZqkaYC
mWkN6BXAykuaJYDDC7TUqQDhIhHXg3pA7H/9Kgf3W0lEvOZyy1VtgZtDR6NjPbV5L6kb8A+x/syb
qHErATp0Mn5uje5Za3bh8ikvUnK9nKp65gd2R5YUJaE5k4Tp0q/bxps4byRDvRvM4c7hILC3Tzt9
acf172RF/3vu7ih0VKW9mBjzHfzBvoSxNhoXBPaZpYxCTNy2yfO9+ZdNt/97/ZiW/66h7iaYnjAu
OK2UtlI+eCG72MzHPkD3i23ZQF02TLyNdgoEGlllo3pDwuj9w7vHFHuzabOMARrz9PNESNsmglss
7i7KrcsD6JTx2hulYkJqKtG0FTLDYeZdjpee2d7VXMkfmDy+n9MvuuPd5rFGsQMMz9yZkQmByafN
dLao4vkSRrq45W6yPbLWzkfoduOqdU+jvU3SaJbC4D+KGrt/LIqy/LiMbPc4vEOAxVhSFyEMNB8+
tlNLp2wG4eqbcvLG3lVED0lHFNHqBZvPZC4OrpaFiduQPGVJD4+3dB5/UuGOYyqHaGzexa6ZbD8o
a5+koD9XgA5tT/s+zBNJzPzZr4ynM4tHOZmbeBBUrY8WKO8ottB6sXX1vStl+zcOGtJyhpFO/ktZ
eE0n6as89FVfgwQH53IhvL/08mk07ua9220CAqDQEZti+Pkm2P5pfFcGb4FVU65TRSn3jAUQkTg1
w1ktJPyUHfGrq2Lx55nwiKl6Kf+awdv0dt5RN3DT5YuZ6ZoiZVcaWwRCAAypV4GFZT5UdOqJgkPn
PjbwQYpoEIOM8AA6mldKEfEhoIWYaCtmXP5hCAXPpDkGiPH6aEIkNOqNr5KH/yvlStyQDvN3EySb
TJxqwJmMpnIKSqZlUVocE+HhSLLCEuzxSGKg0jX9O+wRO4Yhd9NfaY2YtybI2K+1AUpyrv86T1AG
xqIK4EZ7jOHfKIo4P//LMRxLnJuup/cOJGnVg17nSObLiWD5jCtg4sODsbgKsWxIwhNKeMz1EWja
MvdEaUq8/ToWMXpmDDDYfaJfa17+ZjdBoDfzTkEIHIsr7ivyVc4pj7FoT6UguZkifq4dJqom81Td
OvW8lFWW0y93DpleYSa5OZliCrFF4Cu0JeP6YmKntjp4nB/2U6kn6WO3p+n9WO5bc1d5FVFrWVD8
9QM0Et47rrc+hL/RQhoME8Mewh2zncR3D88wb/EQFkF2l2twZgQJxewvH/pXA35JPTntcXG9+xR8
MuhYqw2y4Mt4As98BRgWj9N0lMMGxf9MdOhnRWJQrbCDS3PkZEY3cwXAtN9HV0nIstrWHEegk03d
9XPA5gR8IAFCPUt2N1f1E7vRBXtvfZk0SGAB/RfoYR/a/+keLK9GfLxfsemRcqn+03fb2TEk1lx6
cK/ISzemPrkZpYuCL8LlHlqsxFssf6ZnUTpOgJS1FxYjNP3o9iT/lH/gfIGLg6i8R59DY8r2iiBT
cLlUDCa3eP9AiigsiSREMi9vYaEQoXlBzQelwbmyqg74ZjGLMSpY2ijuMhZ1knVDwssYh8eA5qE0
TuDZHZIREGsNtkfMdPAGpyYF1HE+C6I9/ie79Awz26h55xCEV/jjwQM0bfDbzKfMaXmyDUca1+AD
Xv0YUwHKRP0u9BoHXRu/M3o4Z0y5GNw3s+qvtIl3vCgZ/VsnO1deuA7gk8fqPXbSUApJXBJj4NIc
tmmBpnOmIa7hcLlHWWwnrpcrqOH2ZGLAcN2KPnn/APqRGpYsSdneJialVyeqgWUUe7yWrdBcxuwu
Wl4PsSt+cslL5q1jMiPB5exFCR0NYtgLlQMtMT570vVTXkJxPkxxRbAU8C+OehPWdW7JD4pjZi50
ZKYAPBSpEn57Qe2Ce4IblqK5wB4VktFVc5B00ncw9EWtL8FNeyYvRs+extmRXDo9vKe+5GI5gcKv
P+b1RrPj7d35Uw+UdvdSdpfpbssZWQNL1F+oTXACrLuNwaguAekHnMRYHT+PUr1OVzrrbAc3o6DO
5GneDsJRpaKe0T663vXhM8VVO0lrJPE9dmtihfoIm1U03q7Jb0ksFPjVzKVCxcZPMmJDp/yyEJz+
OC+hdLDvH45Yl3qQYU3WsW/plNfX923oXIzG5rRHIjtECH10ESWutWGr9EeGgw2DQjkLI9cegCUT
W1/Al92e/0OJ8h/qvjJDZ+A5LTK452d/mI8y01fzxwNi4U8aGi70ADHef8qm63bBb772Bc85+Ccx
tcboC1tnSU1w21WACKB5ptpuBLlZYjtxPA+Va9VUIRZFSQQe05NaPlNdtgLlujz/Vk3ktHSaI5IR
efEGwSEqsPAO82aHjyoGd9t+ANjShlnWnVJ31K4hOcWaOPqrlhrVjwC+GsgXZmwyulnnFVZOiSZk
/YGvhdLG3nCJ6Lpcu356brTP4hLP6Sdw2YO9hCgGmWdfH7LgVXCY0kiDdXOUsz3L68Hvd1aszUtB
1TbmheFMI25RxW4seWwVQNLH99ANokHO+D3nTOonsC3VepYCaRd5TUAt16JXy9tRP4aX60oZI+Vd
Ef6n3/uGKmMecAlKz0+oHWrsbB/XdAKauDLcJunWKUHX7ek66ZNixMmNX77xl0IbWwi4PPT1yUnB
Pqt4Rse93ZSEceMW09YYLC8flGsV31KYW7E7jBgBO96Vmp0Vz4UM38+y6QdfufCnkKUhZgwq6ZGY
PIuWCSPLdj8EyHaLNpqQ8n2gw3wpoJvKUewyz3/YMF/NDNdeAROWxQlWjxqgK63l1FE35zL/dogc
/8zMVAMibFFqBaUpjZ/twM7eq53+nfILvLQhaix/X88naKi+timlxWKEGYTmTtoKzbhi+CoHdHu6
k3damN32FUzLTXYC7DwOaYpu0YBLE53WCHhM8qEL4VFAWXY/ts6LMxWgzmOvsE9Qq77wbdk7sGJM
2lkmBhNNz4DGJuRDNkPBoV9yW8I7GYM7PfkVAU2y/QVOeeOc1YI55sJoazwzc7P4/5WAJXgkpARU
h+tuz7t/5yO1s5dbVuJ8r2TPAqmVfBPM0iJZDzme6RXqBl25HtGYHkGOsGonR+RxbEqtFVXehk9k
zRqb3T7kgynaTH8XrMUITV8vo9eSl3LXah4QqWnJkRMb2kk+cVQNpqyrDXa+7tqYup4DvTtr1Crb
6QUB5sg7xIR/2yrmt06JK7OQwGoMAQiHgeMI8O1GlxMgdfclLET23vP6qYSYlHgiIWfiqsHfveJ+
AYmOt6K2mOsrIFW6RazhtUKJiFz55nc3pBlYurTfmS4itPPnWcTW87EHkT+nC2mO1LuvgBEKCN/m
EYCflRnuRE2H2uU0rZa847d3z/ck9y7gyrzGyqJlLr09otMVZSGCVRKrq7gsIZJ2LdYbQfTIneeG
uARfNklO7kfH91I9RQfJpm9/OIJZ7rpYIqVS8bQSZacr12eyzAFjEoLTHapV9udRTaN0CMgKR2qW
sfq+a+kc8cnwp2XDNTQFsGrprZ6w4rLLqdhlcIyrnXhnOmPBuO7vkBMYs9xbU9SZEplK8ozKZHw6
P2+ViGm5cw4/eZBF04oEI9auzForg4wBEl3X/GGWVexrm5QRKfP0sF+wQ5JqhbrLaONFLnJyu3K4
7wxRlrMuo4xlNqMLhBPsf+KQvXByWEiYkB4XOym2iEZaX7L4HlZ5aVkkqIFPB+P6q7/Awj5PhSSw
y3Un/499cDeztioN52SConBP7N5MZlIVcNXIi83fzWQcwl12SeZzuRvhw4GuV/VbkZ4+h/Psa0TJ
bLUkALMKGt9scMAxkU9X5afXotPrFhgg3OKpd87kkhWCrjZiVJwQESfz6Iku+69+FcAmd7JWOnDF
CV/hw3Fs6pW7/YCQDtCOJV+IO/SnfN+EzW7vgFIRd15gQ+tu/fP4l5//T/j3fFbq1qBBafarOqVl
UZaqoSj8HyLs535aRkXGbqCsuN3BbV0jsXGfH6o8HJOc5gog8W/167IHnHrDVBYJXNuncJ6uhghP
JOHWrRhj4xW4fjUcsg5fo9s5ZzLjoIOxi8fMNMdn8IC2mVaRLKungxqFMvC86UcwRGO1Z2QcTyCl
iqOmR9bDs/j3o9PtMiRafOK98Rtblabtdr/0sk4dZ8SmfLT0jmlHtv/pbh04PD0IY7N22yvrhyVI
nZD/EXJn8nXxISfbSsRg+xg4M33S4EabiVMCD9Fe3VZpeZH0wWAdvMutdjZKxJ2ADY6rfKbz0Q7o
YImM8NPqklUiNRUQ5UEIESnyegBpW46mrwa7mPP2APehTgO9Oe0c9yWcyoaOWnjnH58GQvp173ii
zzt/pmDEXqdGV2kQ1d50XgmEBUwk8S0JL6KxqQVR6ArUrVszs9+NgjJWVaKB/oqkkmbmgzLXCsrb
25dK2qswjFz8035FeUQhWIFvbVLiW3yfxrgFYsd8mQsK1uQqT8FJ+wWOa11zG/nuXayvJwnIoEif
A698UtxocqFQyz0LeW4um9R3k+j2dSENnkWBdJ+ZNO2u1b75z2YfmUzI1QDd6QTEmjOh2B1GshFo
z4Q1MttQ2B4FyGdgOqtlA0hEhRwCtOOae7VSafoGi6BUHPgXos07x643+eeL/NFpOQ0sqF+kTqvP
2swsjuGP4PWbPJoMH4lRHa6UhtwIv4wP9xit/mBXTKxOru1wIqqKd3wI70CejrfvoIu8IXSpzf9Y
GSMddq5jxVrpXr1C3IBmMm+WqpgYfa0EQcy5NbnIp28G1qCvE76a1F7eoQoN/mhZpwNo//mOUINu
QIlUn+R6SKyhktLNFeWhygSqSe1qwMM7hIoPMg3lZNLIZs3DMQ4mUEdSSOgP/aQYIfN7i7As2wNk
wdQHpmJoYxWvNPu+V6Ku88eQq9oduF0uyCvBHwOc7pSII3UrsVrk9RhdCTT/IY9PWdnCp5l/63to
PSM3C9XygE/8U0CYnoT4wyl/SGlMzfltVPJmF6yjDl3DyRXsFFa4shsgn6FBpOvqKFShvKzkHqaf
DE7vpzGsv1AfiE0xaV4W4FosthL5HVVJwX24EDNlWiqJRYotHknU/PpES3g2sl6HoiQjtR0H0nP4
bCLkLgZeSC3kBy8/Co0gTgo7ZtOd/oFZ64INlwg/5hRw4cqgA9p+Qv4nBKtpbWk3xFyKX9b+b8C8
pa4areuXx900jljN7TB/8zCNEa4tG/ogFjZqD4Jj1EQb2QuOehGbHtUuEWPXEQGCrRb3/RN8ujhN
qLdBZg/Jip109cUSj3C6JC3VLq+BRyd/AFNSULu4htLmNYpBbX3E1wkhRuW4HvRLPZafmLZsqXIQ
jwjOWiYXQr+hxV3Zi0tfQRxnGGTZJ4pw1qdH0DrgN1JUlfcssW1oALoWNesj4zgwZyvvta18ZRSw
XHrbVJDNPsHs38It4qlWHEqatmJ4aKR6Bay1lrv1XElU1NiP/AySVeONRFWwOOqJMVxaIAnBi64S
TqMD7SyS7p8cV8jx8OZuKWX9IkzNF0dKGTbB3iT0pPuq/UBoUww/mMeY7qRCvmBs9HoCrOnrMjDv
D8rWfU1A+/2Z7ENU0vMBphOno0roh43X0JopIUARIIAfGt4dfB51S2PsCPh12/RUch6pTZeZkiwq
OhKWtUQ7Mdwk5ngfJ97qJHv40q2tNThjKXs0b/DpbsUKUpX2Yeer/fxMbKApwEMOC5J/ulv7FaqK
Vxd2E7FLX6PL6HIP6KPtUohQguP5OZRiIcCiuQQpKA337PVa3+W7mTTs5TRzi9u1aDHBsBQQSXXQ
GKheHlZZK6+RHnPw/y7mP1g1h3YvZo/o4fcikbxI9rXimtQWOQDw0A9aFxnW6A3TAvf3Om52XiN3
9+W0s4LbAWlmpnfzqr4/HL0eN0EPcTw2rKspkp5Ip+WqeOP0Z3tqlh1nxl9NZ6QFOLeLzYFHhZfU
TqQGyBs9b9oacKXIOtZUGRxFr8zlj5TD9N+A2XCHyUEDWtmy9u+6/5G92YwpBDlC7eff7oFoW+xE
cPsHHKNIHVx0fvk/3qsTI7D+eXvmEZTn/YiZQdsdN7crl9qg4tHciIKaf6wO6SVmNtyitEXhH9er
AQUMKNTkY7Y36rjGQFJQYZQNUjTwRhJ5/3xUTKNA8wBNIpU+eh4r0iWy1rkB19KENnU7fKisPBcm
jhhIpxk5fDA4ejDX0EIfna+fiVeKNNScj9kq5i9XhczGmQpaKAl8i7oD0XNEX3MsmbUu15oMAMj/
89mUuCnf6EBk1uxxS1SAfSTNYn0liYDA1Q3a0KL5cN9g4kB05vxyN/VOs2n3Mvrz45kf1dI7biZk
czWfUuJiDyGTVD2EcM14W62w2hGrt5IFmUpnd4jcbwINLAZo7YagkfrlXcbS8mBs8yDaOkP9e2IJ
2FQWvDHs1vfzEYHUbwYejro2hXb1OidutEVLTQe0zWYbSrFkPuynLSvH42C00IHYEQ/ehZGPYgAP
1+w24vXHlcg/cO6SbZSDyn6kl2CNeI3ZjyviyyaULjtZwwDYkZA9ojmfj/RiU8RDieJqk1Ev5UVj
tcRV92zC9mn3ub9wcQBYABUoRFnHcxSIq/KsM0SHnsFC6snHfts9ACNQVCWC73BiPyyInlltz9e5
r/Qxaus3PvsCvOt4X6yfQFemvia/rY/P5bFSfuRS07DFFLoI7SdiX8mxoayz3in2pbe5EfJ7oEFK
0iNe1os/yu1teBC6iSlcm/jzNkqM/jwVKNOj32zuwox33LLUbCLZUjlipdiQFp+xJjiVlyGC/1ED
cWvQI3WnYeVx7I1biG/xAvs1jqwgI+n/MAwht2zKorNL2S3ttjfn8yOi0PX7IiVw0fXjwjrNLQaz
hrHKCL3/PJT3LntrMIC7/aTRj6/LBxl5tBpsXNeKMxYDyD3kfYileaoot86FIflVYEXkx5csblCn
wAcanfk7W3Dt1SzIZrIKZj/WwfVCtEnO6U/TxLlNbaZmPYbmKU/EVoaOggskCzoRdFSkWTXez/9+
Z366G/+v5YXj5UxXg+W9PPTxVf6K/PQtCKNfjJGEHVW5yweO2n3GQYrZuu9PJQiXCA0+Hjhpip5W
GA7ve7jhVsFI5fNkU3sCk2niVi2iogkxwQ1jxaXb8i4rpGNTXGMGYbceL4o9ieCQWo3J3ODSZrb7
OXPtbrkG9BOBl/bR1veMc9Kyb/apSSn0pDCqtNxwMMrKZx008IRnOIoYpbE+EB7J1beMJ58PfgHP
TFXLHW3ePJz8RIb+95ad0FCrzQQUwj9BNYO5xGM7fEt/YbiUg5bY+oF02v1CYS8/z7wcK4X4kbh1
F5aQXlLHcs5aaHlJeKExefO5HxzEaA68i9rAgDq8l9bDNHruhtd1sIcP3vFy0/fn7EePbNq0MVMg
CEQ+zQTalKza6jgKcMvp1boThJVq6qKWCVcS/dbxtU1GzbZXwJw/lsYMTPSReZnJU7no73XxC1ol
3qGzAt8wzpIqqUyesr0YyyOtYGVjjqfFfLsSkMFwsfiXF3dxe3PNYZBzBk6sQOpl2FDNxo4SOtgy
mNriDbKl9SyRyAYxvbZmJqNopPfSw6a0DMczv/t3Gi8Mixvd15FarvUWwl5xTAXDapWiSnM6LxkO
3mnXQwjywV7SPG1VWUOLPFKXzlc6gRYSX/ThcT3aOMbO4XOzhTBOh/Jrn1NoP7QclatQHGCreVnK
b+ox85bLuuuZO/UVafRCfnzdcm0A1Hz2ktyBoTU0WTbANQt1dMUUoCEMm63/VW74zFS5/Tc1Yhhv
oGOX7CZT08uebv/Mz9fOTZl7htEG5hDZ0JP9Li7M3qmIgz6C46d8xAsBLP40T7r6cEBU9QzppS3C
PVHWEDu9KMhXrEyvH2CWFsO0MTYRrtW3Bsb7lRK+Tqr4NcmxtZNiBIK8AQh3PRXh1e2sqsKEjcCo
/N/QD1Y7SZ88ChhYe4g/fy1IGH7WUL17X4Wu0838dzr/tqXaWDS3U+9mPB8ynor35k8wIsfRLvXm
JLNaHHjzjb9ef2cq8buivcNlBJyjBf67HC2yzK3q9nGLTQR+2i9GDBo5uYuyhLq/bXQSRbFf2Njh
7Ay9c6xXOcIO2T1jZqAI+R0HjmcXkvgHx7JBZC4Bd1L7VqjJm9ZOMr9ip8G61/coBtiAafpStN4I
kdsPOk5jtAknVZSdEJvd6Uz3DuTasDxJxK6XEp8NtLywNlsFzfmtcDbIyChq4nOjU9EW06LAV1gq
eH9I6sDuyNgFk9T5lzL7h0qbouk2MB4bJR4YoYl5didBLneKVMv3b68AwYqav2RyHL7AwDViZsFv
E2PbSUVgAJNrjrOx3FRmUhyrbnqiiIjT/C3Wewr2BofX7acJqPk+KYIG2BxZE5AoxYYXah7Ep5jx
ihDT3PXDEq3/aj78pNHQ7RUSY9vdPtv19dba8lwXHOdvWzG5RaEBGQssJv5/lFGniAWzUzFuD3Ld
z5ub1GiSsrS7lXPv7bkOptJAeo/S3Zx1HZzLJc/7uRiqpyvNqV+UcDmQ9qscz8pMnUt4TY1jKfDc
XTCVk/nQmI5a573oGgKjYZDd2lWyR289TIPfmSB3y+oc1TVf7fCiJRXKlFwLoIly0iHzIai/GXND
XGbkoH5ee2KBEWBbDFzC4w4bqRWt8qKlBlobVkhoIMSt02BLTtBhKLmo3/Sif+X1y3xC3M7DWI2e
puWk5TH8W8RCbjHxTji+TULpUVC6Zv/yxbXkPcUL7u99l2ywoGKZqUiI91Wv+eydcIOCdA6rpym2
bxlIem4fsPSEhMzvCLuJJFOy9VqPwN8W7WaTtfuBOxE/in4CtTSlDN0dZjoFfaBpwzTJvUYHd9mh
6fLuSktC7U8gtkgP/fiEsMPMPEHEahu+/NI37IXBCAsSdtVw3yzqAXbiG6pIVRZ3TWgTiRQIX/V2
JGC60GfHCJm1a3YcDZcS7HplSZdoU4dvtIOAxhw4/oHLyJbVku1BEbXpT6tTV1RM/v9T1mlRioJv
58pgxfFNl9ld5nBKzfDYTvi0SwAlyLAgjjYgX6KnRt5QGtr6yilx7e5PS5nee/edH8f1LsbNtJ4a
iScYtLkdikRoL4J/uCJSS3B+bjs0LF0pGb6g6HVpo3ep3g8WZ8GhfyMQEwxEmVijUdX30RXpnaza
EtUfs80r9IKtU15kPUPwn8TiVPDAX5KuN5vxTU6WOhtxiyCfdNocnOitCApT+JbSq+0QK9OkBcML
7Hp6a1gYpeAcApqMbMiFd22L7rktVyaWcG3SJB6U6DOh2HXGt3k6x5bgf8TaU0unCLDBot4sc6Mv
8PptPyKF30RwN7KWAVzrRJjBNkvff2jocdZCqBcuYzecC3PnvMY5cnpD8S93m/nrysHjusIiITkg
rKfHZBHlxi4Misdo2mvxIRFjRFOjms4AjkgsEpMkittG3mAw51kmEidBtRLjPO6V6YMED3RkLv7i
vYp/PCExoYHyDAgIXjy8VfarQWzO5oQurA9KT8qgauCaPvEPjRz0uhV32mJR0H7A7SV+3SJgDtaJ
4WEHNVCG4XXbyO+Ks9p2qJ5mBY/fS9qs7vgK2qvzsbfsX728gjvMnGvNTMNi+OGJM42SdYMXhZBB
kjdvtlQp/ZMrnkjGJUX3EW+5AGAz4peloymQmYeR8LRiHgg9rtkiS7vd7odzuSkmd+5o1Wfpo5OV
CjEqvpbCaQ4QM49Qw42KvxjX8dWPgeqzUWt9U6K427WEo4imv/qcbdkYRcM7OYFr+39v/rhAnipD
0lwFvYh5Uz8qQaH5dc7jkA4DGcJNYZ0qnN6qP7a6XFyJWxtzH2Rl0f1C8HDCCC8NouV3Vk1/oLzN
DZtTKbK8DsVsFT7ituq0nqqkm3WEXMfk4U7cw8zjexj9+xG1P+DfM7fQzP4NjfwgNX3aYve6kHKk
xXklaNPFinQjgsDcfnUornAPniEbx7GdXwG+iCbwqSEPyuaqdcewGCLjRpdm4KS4R+Pu6u12Q5B+
42ZAJ5fELMLHotz8O4UxQlI3RQ5+Hh/PGCfLDjIEZPksHhiEmCsjWEj8UVwFN8ANthdwqfc/dleY
C1yVLEyisP7mi03NGMI3K0RBfy1vT3OZ+T9vYOeZDFHKBNIVXpXs+cDqa7IRTiwmv6+oKd3jxxsb
qDyH4li5AKjQPb0jKYzbSaVH5dB6qWtwpcO6nprW09ycvg8Pzp5ll33g8DerWgVRGjs8M3BPoLDG
54PH6Xs8s6OFnRAN12S3hvD3lEoOokCOD8cB0zZ61M3vvdvGz3iqqZW14LwuJmmK4EfRLVNthik7
RIbdP2GZ1nPI4hgOqLr/9qrUZRIk0tsXztZzUgbahz1OSj1DitQwc1FwOtMlh6PI1XMkvU2dlNpd
N6QNCIl9GpRCUds2502gB09aEU0oHnAMOPcYylo6O+F8WwDGMZucf5D5I9EgGbYUEzEQW/k1Tcp+
Z9xPKWSCJwX8EcHNA/Pgr5UqkCJTk+IIWPtQQVh3zA0uTFWOq7bdoqUzIIBM9BrsLRQdesbAvwrd
rVw0Jor5unlwj1/V9ZUmgeCppRdbpHJgVNsGaBkiRsiJIZrErd+L8r8elVzyw1BJDh3+mTj++TNo
sJBenBOaBxFoLzh+OBYPLsgibPAJ8bcvyUdFI2hyYdcPnBTAZpXWUcveBYdXV1s3r/u5FvHynm+1
raZM6oMjBsYSAaeb2isoUEFeGeLRN4t6jZSXtPFzu75rrFG3I6hLHQVsWo8S61kLTo/uSdQBbm8t
yZLm6TgZHtDxZ91owXq49k3rKZq2Zi9+YXluXJG6INbyWeODpZcP6cZhJHsj6kaLYjPCVxvKE6tC
sSzbEXVrfCXRF/+fp1ek0zT4+40VnFe+xhykyF+e0N+wA0x4bDtOXDY/OWbtIfggJ1WT6MNWFGio
n9D1UyWuhVVV6pqT7+EDFO4awoC/j5XO3gtnHy7ZKosJDSBVgb6GDGygXVFncA+emkevq1pQHWnP
jD6+1i6XNxhuGf0FTVIPdH+bO0L59/robaJA2DsvXknJNeBOvFlGf1s7WCHk46kBWUdMFbbPeSLE
7xtULv1mHyRzMJcrkI9tmBW9uEOPx6V6XugdIx3i4PhswulM56mkuinDuOZCBwCxdqCBmLlVLYm9
hC7foi8KkQpY2FeCpjrMhjRNuuThHn+jJKnWMuSpgZdIz0NH9TMVAB39heR17gT3/alLeePJzUT4
ha7qtZpQ2bMTKzFsx0UnJcvH+2cvR7IQK5B7Yh5PzwilyA0T3nk1NVuKY/Nq0FlZI3NoSAtuMzM0
RHM62/5t6BDs4KoV58NE7NChAsgfPsXIKHcCiU9ewZQjOL3XC1RD/9WIpnTX26FC1PE+GlerR5L4
1FBkvoHChuR9phUPjT8u/RRFHsT3qre15BHXsiR/34Qd0sj3WJxip1mbpe6f9Y/1op2S69D5CkN4
cQgnM4fyf9dpR/UVNighcXBH31ldcXIkLoMFiWNJBXd7Bz/uJjfVsSkyL55uiukqt8aUxsJrEQAK
tkiwDH6giYeVQet4UuMjgqFfmLPVNxqfp605eriIzPrCRBIMpMPAZh00aJtXYgHTKX30qhzDrjSd
EDiVFZGn29JvrMMx0Y5iyIuSNVjSrF4QzokIArxZD5W7MsBPh6EpHmbZlUuK7eijvDtpsZe041fW
P8qEebYPElS6znnU8pLycwg969wsqAVRDyL+sHHMSXnN2OHn+fX0UkdsR1lhUhZtGhnJzchlkKa1
a+8poUz6piKtyYmhPsAKZtO4v4zs1SHbeOHBmGMbdXVDCTE26fzXMoc1583CruCHqR4Evsq8Y1vf
BEj6/NrrUdb/TL1hgTt6XB1RVV2W++xmReVu7ehECLc03bNx5BL3jPOu9d4CE6k3y/pB+fd56Skj
QbTlveUUz2a/I0KH6qbYQ5/zNNqPrqFu/ZjC4/gvwQCrYvPhWaLY6p7KwVps4pfUTp/XrAxCovBe
2rD8TA5OeL8s9tUTHVWcWsUi3wXzDmrShvpnWIilea8lm6J9d5mvzCwiMO0wX/NOamCtPBP0qzYR
dpOyHVswc5Ixdv6ej5jkkykUjtHSPYE2MK8GZ2fA0URfHfAmi4ur+WMW0WBdZWxbD/DsWm4Q0v0n
vxTt2Tv8bsX8HTenuF2+ze1dZAGkffVHgAWss5hpT0rks5TJGNle6Vxgli+LVLOhVKKxLwe/rm/w
7+9PzejkT5CWQ+CWBbvcRq+fq/utcA+/hmyBHJgzN50a1pIFv/v0FzX4Gw5zkwOX1YJFDPj4uyP8
tarUIBArhEwK4PJCsUeiy46gQGRujHcSE7piNrbQOmmQPWxqF0Co66EZS3E41OcSV/as1tgs/wY6
VFlTU9bPsEEngLvoWH5AeETo/NETnxpA7fsOcnS0rHDHVQbWohAWWdXgoJeZPqvHd8R2eAVjtbh7
9RTTS+BAdrLB4pyS8UK+90RcboK25Kz5mpEYM5e0fNFxVBtYfTVZyJLwwOleEcPnWC1cKNYya0tr
AQT15rQu2AwIUgHrRyUNx2NmohRMDQBL7nvOUqo0kam4oIc23EaPyuKT/8alHzSXwsLZgxpdbRHf
tjdOWSewctHOGoUg/a0j+u1ReSgaKHRQ1NlAbf1JTjyS1knbtUiprsAUe1moSw1ljn/PWw+S6yZF
nfuCJcLWzhWLULd8ehzCpRDwA+29VmRAyKz7rm7HnPxbEMQpCvp6uJP4KYuvw1h1Nyea/QgyfyNo
9mc7DXrrX1WLM1chMNMJp2/0jHR9WIQ6R1qIhm3chhJROs4vKtFaWlqbU81LJU6aEkrEHGSkitzd
Az3Uk30RGd5nN84UDikgHvd6GIBQ1xus0qKM/Kz4VpFNnlYHjH1y5mIwb6MYICTb5hvYa+QItxCP
5iQCvWdPYXXFuEBarrfGCyCA1mJroGu2i8hwHS0f71YibJiP5FGObBhrtp+GJ0cQiDX1YoD/6xlI
u3WBvpccyNqq1a3biLaT+VpfZLETpsS/rYWEgHf9M5yAIXcVyJ32XznVenEkOD+UuyG1Iblt4Igf
1liPazaDke2cQANjHIl5+Q82/AImj4S1g50ON/wYFfYuzwr8hf9llDeBRXp5Ucp87JITlFCm6kFc
cqff/D1qIkODw5zy352PH8eKvL/f0oFNUAkAOEq9/5LHRndqWAAXpKSZY5XVXp7MIjJCwp5WDkfT
36zVjPuZimCuQvO7BSXM9z1ZylqSu5oJpWQzYDuHlsT0K0A/pt6UjYce/LWqyG3b6oufZBwIu6s1
cxe5dS3M2Qteh3oORShwF3lnjcI+6nOi5uSGEhiEfQW7gXBfH1d60O6mAIZeuLp2XFVnP39oDzBI
hT7MOIyJePG3I18gW8AGrRhkljp9T++Nw/k3sB8hYqvIGR7ItiKZRlfHx0ZBifrMyDxkV1Vb17Ke
0KCTGMfcC74ByH0/o8vA6Aj5VK5eyK9IayYfBiXD4FtkMSjdZaRz1L+IJTezQSO4eqxVYnAhEy03
hP5aZrLj3TmHCk/3VgwTwbNmCWzOJByu+9wJg6vBJWhMBTUiMwdDzp849VTmQS6Mr7mwnNl9JnzO
lyvl1ODrSflaneJwZys9yT5PoVyUAtogecH3oEzSsJxcOkafBxPaYLp34jXAilpbNgci+jXag1Qf
pArlYnvfl99gj1CeKpa4Q99HZZUnLTDs1rw+Pf53x2xnLBSL+iurpa6+u3p8g1BuRIevV7ITTck5
KuTVd/6+rD/7iRNFNrXN1z4BpNGIVBOnlwjuomCmVm3522avw3svEnMdxEJjYRc/pQPMbKmmI/S3
3C5YM8yshW9/mFvtV8OLAzMRMXfv3Z4wxKBCuSzdrCEIgS5BhZVPmhwQqOZzkwAPsVxYwA6bqfnR
mgXL14Uu4qmeiLHR1vxMnJ07qHkTUuBJV2aQkAC3dl9TkjT9pJ7zO+Xd5mFa1s6zgcIJ6tNZ2aVr
li8E0VLHtYNNkOsuI56o7PwHgsZff98cqFgLjvLNfchKC+NMOuEnYtko80yo7UqnF6Y3KjHMay4b
amzuQfJNo0mhGqnjolKtrlJtBcmVaDmgLb+9nYqy6nTgG6Qz8lgNcve4uPMw+ar+vmL9+hgUTFop
C24peK8ITzWdyNWch+fkyJ272ppEJFEAUT58+WB6/TQIZ8CUailo6+nyiiRMG7m0ekNrk7dIak3L
bxeB6KKR+MmVSwd9f4cr7jNhKzgIO7eEBqPfqVwBZ0YnrVUXQkxHAVcoFUtlrZ3xzKLr3TN9nES7
qNxLnO6Sgj+W0FlszJ4sBm8C35/dE7G2/q8n4xqlfv6g/QEv1E7nypAMQdLrMBgbIVxba3McZZsU
aoPejhr3N0KGY1aAzRMjAFrWNhjQnoYnk6kXeFd3Le7LOlu4OJdZ3AoYd8mpqOMkuXAuOeo31jxA
mOdPSdnm23E/RCeuNxsMJxIoL9wfWudvEpcL0UuaWtB+/0JfXbreK3r6raiai6ckK2kcXpzei7jz
3iCflygJzSDkkSoKLbwOwh0haTtj1KzrQyL6NWqVu/uUwcQLsYbyLHqEgf5mXRvISyVl0gCI9E6e
nMzd0+2drz82wzpR/Sk6PReuZYKLL0IIM5IvzJvTMdKVrutCkNcFeh5C300jywCXDfJAZvLAbv03
/EuYu2RCeHNyYhBfn0a2G7aVIF6wzoN1zi24hpljxSR9vH+3zjdm4lxo8H5XP6DBhRpxu2haukmF
ELyAMxCuBj9fSazOUvTsuxzmOtMKHl+hW2D2wbhcWc6TUZwFXdch2l5w3rjN+xY/O687lZpZRT3v
1qQEnJWzkOIEGyqzXjsjCp7DUxZ1I4Qnr6wWBZoYrAjXZyuPEKutAky8qEeG1Gd42SjDt6FVRJ5f
K3n/OQTIN/Wk+iUbfmdqSmCZG05EorMLhBdwxFwq8cpIH1V7AbJbHaF6GlYI0qkGRA73q/pwd5BJ
lDsU97+EvfO+31fkPIW3LxzpxdsgA8Puhxhxldv41SO1/wstSTNyYiKvXvva7HnbRl0dJlrnsBOi
2qK2JRtsbDqmT9T6DMENxSG+kGrAOkzvEgt0Y7hN5hziVBbo0zTsmPxsdVhv/7pEBghywMKL9cAs
kqbhCg6PoGpfnAR0unLCbfvL1Ah1O9+AZqNI5GlwyIMuvkWbXypbw3Wt9Db/n4+Ccy67w9yIhxji
kDYj4gXt8AmL6gfOD6gsROCo4XAvi/TQy8GmXmlH37f+fEE91x21BY/WXWqB2Np6KdbK4bq5v/f1
kZdbPqh0LFwcAQ0rlJk660UwX09C9C6r2STSgBUXRCaF2jPOl0AlfUu9BIgP7JlNmP0xpaFmIIYB
tqjbrd4cmmzeu/r5q1yXzP2A5ZrR1JD0r5Irv1v8W+Qas0MRAluwHMfXp/AW/MFuIw2vmvz1A+0J
wqPfGdP2q2ALuU0Jwyhbexlj5U5xjVO5tdsLMXYCK1g9F3bvfTNd4cK2YCUQZ0ySM9e0844q+Sc/
moWCZYrEduZJt6/qGAM725F+58GemakUMJ7kVcep9T6QsqrMbSOtEoJ7fTrYHABVYHjHpu7qnVsf
l+aZKzGyA32w/nAp8lM6+fHV0NXn7wp9CAdDdjfw5ysw+tN+SkudvfD+xZJyqU++BfAteUWPfFwm
SusZ1EMTl8G7q1WQg9g+0uMM35MIcwBRMTbctFFiu4tGXIXQKsx2sv2jxIUGQEQCll3Rse6qwYG4
y2Kh3BcoGLT0O1K7qmX1XbrPT/E1uo64FFom/0FN+z+/UITMlvLKbiqNsxKM3KdxthfFJi830Xut
50iO22THQacQV8Ai5sc7hOt3UkUhsu/4QHb2GVYuRR8SD3kQOu9TL7+r+b48czTVhJ1KMJyA27qQ
fdMlILN1YIOjgmTv820Vz4Dbwn9d2IwzxCpGG7y8jRdVvTCy3C+hbrqIBZdDab6Ys8+K+ZeCXK1j
4lEJdKq+3r+VITqok/l8CqL3vIemp5zeMZjyk8+MMAjyPnt1S3fN/a7yX8/K22FmCymG0qPH8k7k
sLISlg6411SbJJdem9fMufHp+2R4P4A1Bx9enPGBi9gDlcDaWJDdvqTd2kWipeHbjwpa/9xYglli
F+/aV5yqh14KKqEpoliIsIzvCM8Eg7mZvvwPfsdwK0aZDcrFIwaZud0OxBiPAQyBnXrbXYbv9HEG
g+YkPJtdEawSoQlpOe7iUnwClJH9jNdOr8oqXDQ1I++GjaLbhPYSK6/G+zerrUC8hCVUnjG0JGRg
hS4d01/Texuo0EMvPPPjjuL5DQN5Az8PykhQxZiXBEy8xV317Lvxt6TqLdvzOvbo6nworsWXi1lp
uUMY2ufHmqJ53+JEMDGuE1K8Z0goekLnZZd+dKOyP8Y0Vgeqb1TgQLaBnCOzpR/7HOAL/1rrX9Xd
fhpmZnFne4I8GYxC7y2JRPc/98XQFxy5fUf1l9KOEwKZWARwpUFTPF4niPQkZ1mHnq2Hq8T/fZUe
Ce+CVRUQO9sGGKjpsNa8h/kVYbUSfb9yhxd2bwYkQPpCAC1bGZFmelDlxONnWGensjimB1EvsTZq
Jq+nIyqUUTPyoPSOFtpB1KPmNiXEcYw9OkGOnZ4JoH2nCXBuPiOZA2KTfH6iUCOiN0PpEsIJPr/p
Q4vht0rIqwWFaoIiTG+44mdCIeHxODWHayeoaeCzGHgTfCH6bIzZujOFtVEcNn5jWzmzcQ86c6eC
ZFcG9IPXrJIG7j8r7TnywCEBSbzjwaoaEu/zZmNwQRykSsfV9oj4XS9baxSZGC/3F6vZ1ONBunKr
Rvs+rdhpzjPbZ3xtbTDFnsjDomFOoZDZ7wcSSGLm8FoxWQ8k5M8jzfxm80Fl2/RhvZMeZ0yWiu2h
2fv9B4+EuhH2aQhqYyWL7fcuj0EmcDgX5Or/nMBvYoZ6prqFjURFsu7QCIwRGz3756ZWHQUjw/pp
y1ywY74y/5DHo7Xacbycd3jmeDr1juT9eYRD+X+qo7HNLgHyroX1+r4LW22xm1enSfW44GlpAXOW
Wepzv5rmRV5Lm2y5rm9ptnXGahCHJaUFoz5LLMz19cCUf+wp+Zj6+3WL16evs7mplmFclE5+nAD5
uRikNFCawRb8qu4yQxa1K+O4mT4qd70OwpxZ/5SVBUyY0aumozrQGMBiZ0bcP0JSGPFXyQAvd7Uv
0I8mYJCJvNQnqJ6He3Adbz3FJhWHDT0XspZ7AmPKSh4XXRYq+oYTTVoy5hxJatBIsma6BUPOenCP
tW0N4W5QKhnKOhiNrSUHbcTYPgNurPFtvuEuSHsoIx9tH5/JXuS+OuuSBUsNlub7WGUypDMMDet8
SyoLX1Kqrwt+TPM7MHg1AogpaGcM1urwrsh3uUHICGbLGhVvjKgLf5RYoMuGjh3zJ3Kut0UMzpUt
vnUNn/PoeeFvR+NQ3iVnSyOzNgovUbWsZ2XMjTw9pQ2MgpaoEdwJ8gK4yH2VxJXdynJbruGdSOxG
zvtFvZkT5GN7o4SsgTeku7GR2HiELoHWVzbGsq89tfwSqtvoNXsUabUaLBrFVpBwlCV0/SZXmxIf
NlYtnwlv56KjcjkX/fMlOb/W4Bssgg/xoIH7L1BH2qg6jHWBr2yhI9l9n639MFgAUYZM0onrcdcu
pdztIJ5+F6mEjQRTSNGD2Iu1GnZnPP5hyeTslCRhBtl3S1cUvM1IuhfYD/Vjl3P8BTWZWmghJnag
7pGZj9LPsKdm+BPVtgCEIxNZavEBiqmodKvsYlzHYm7tik+XRMAgDHszVkj1TRlIZxu5bRS8jkhx
KI9yyXyAyofVwdc9apduU1Px1WfeYqAzMmFITE3Z0PfYDx6sR6gjr6/9fxRXfD8cX33IKPojbHCl
YeyOYY4p4ksQ8/Kdby9W+MwL6e5R1fmByOgp4jdrIwp+GYKJB+zIe/2g8MRWwnYqRk+zrROwGZ+0
tzr4UBi5+uhrokcEmDHmc0hzTg18kQDhLe9LvEt3I6gFsX9EIEmBRPXTEunD3P7xMLiuHI0qZGtV
cwnMATnQzETv3Q9BpG+aH0lyqjzlHN3puHtPqFVCqgFNhLc6Vlg+020u1NPDIQVPoqS6+HICZtjm
qyG5X//y717nNvQRzmR2Zuktz3FFvqOOsjae+7e+HjdGKpYoUZaT+20U/lA4AUG8/kc/mQpdGjuw
pf3OLOa12tidwyjy+tTvoashg8mWdS64kgEEl64cd+31xYCkD3UIu9yaeInlMgjXRUPBOFoiQwWP
8U7GjITkIu3LuwrIpWzIDOSp1qBAGfmcnLA8ekPnMEKvdtGGX9g5wHoTlu/D81NpnEvClV6F3fdO
V5QOCLLjAVG4MwpI4I0EcfYiJscZsnRC02UK6pxsFpEg0KoYN6aSPsNHxl5/mtuCvdNcgvGh+xXC
baNch/4+3VaMPc2xbWqH9oQOOXFcXw/maKyMra5ZIbuqSQp2PCBmEK9HQiTt+jLxv4/nWYbYd0xL
OtjuK9F4UX4JjwWaVAWNTqzIqIvBteM3k0Tfjkt53Jjo5aunaC26UVYOmOIg7DQ1KBdLxos91UAe
gJc96zMMDTsR3w4t/SKz1g+w/OEXGIqoMmul78x20h6W4pwYs9Q27lCnV4j5NRdQN8g7vWXEsbyq
9/pVDj/il8m8T7RTzF2uQOH2JQeA0g7TfkzWltEtAv+RhUg8bSzX22Di5lfIF4fMiaBPrt7EAbmK
suO4GA2j4LhXuJeQd2k28g16je1JgHxhhsa3lswAulcraGT8CXmub8Yu02g/HERV+wiTzP6Yhu+A
l4lOkuJMucYizYkl5CLfTSN4iVYAR6LQ91MwIA88O03G3YhpUd+ZMeoY+FFVdpTrF4UkobsCUFGC
xdoWWv2KzAQbkgbR+Clqp3McFYMxsUyoH13iGXyxD9eDuKLt5MJGMcoSry2miVpCAycLsPZa6c6W
Vm9HpRMNDMYhxSx+NUpzOVm6hhDyi6+XjLF2tfquWHLl2D48E54k6y1Xg/dNuG6t55/N1eDEzbay
y0I7LWIEpVSYvHZpKXu8mzagg/FkBtySQn8wn6D+zajix2jVk/eg5KQbFOGYsbhUnx34OdvdmHuQ
CKqSU8u7wHzPuBKUUhwg1A97BORylsK1FiSl5tKPvmXzZXmqHLMooPuqZGzpX0Qqr3GuYN1Ak8xo
Mq1tWxfu+Lidwik4oAyCS7P5v25Wzrssi7ufE1dh20KOdwZBbEeVS1SMTzhspQ0GFgB4oAO1FNzv
JgmtNe+IhSYWKVPSwO9KmfzCIbPCKI98NzA1FYTR+A3RkUKJRSZTgSNusGI+B+75MLaUrr8C5IlT
o/oCRPbMAkPKH/T76YcGW5aZZgcv6+tQ3H7sw5wOrAm76nFGja5GCyLUIP6whM8EwlCP6NXUZYkQ
oErMkvT3MUOQzXMNrIn3WkYvacUANkbe53vxDpaDLv5KuFGWhbM84afHs262whbUZZeo2pUOFxY/
QBMkA0n9kitDqKILC5jcmssfpVm4HOEi8j82CXrrWVvz8fUXySV2QM21pL+F/o46ETIbHevyHAbG
4qRdVzykYsCeZZOT/Db80VGgLA/P9E8VYJB5zRBpbsGRkv2dP6ZfeqdWT4OB9Mt7Uv5Zdn5/4LCN
9yWMGrVRIWhplXP/CJGBD27/baMNV7AcORPhj4RAXp0HaGYTFu7GSCs3heLVXhke3xeVU0vvO2xA
w9BCiE0jCm6P4DKyQf1r0owIxex4Hka8FS/6gTyHhZ1tjPuZkl7v6Em2xOU8sfPCth7j3ZnO/FKS
zsDHwu7/s0byggqY4xaCLw52yIioGSqqBkBsffwBsdl8iuyHPNuojZE8GvmScKMhqyCKCz1fRJOB
PzzUfo9CLUNwiSTCCeTGz6ZLcQXpAc3jBy5fbwKDPqklgXT46b0mHGQ8wx7RUee2lU5rzKC1uTMB
CVwxb6BnoBZO/KOkMtqSPf0tgliwXu7faywbsqFMw5qkouOPQsZthqPPb/TY4Y4NeqQ5dA1OEMUJ
hDSTxqsJJdVke2vct3JSNfxXFftlaF5y+Bv+GjH06VwAtUyo+8rI6Xs+qOAC3CjzK7pw53JswzgS
CW3nLn3w9mBHqa6sDHsDsqJU4gVoLxCXMZaEuq9UYKdXXWyRS6fJfLLHU9wsi2VTUtvDW8m5w48g
671HVP0fQzgy86zkJfJMmEQ4eLasjt8k0eEsTJArXzqT5ypsmJQgCMWn+Hnlm/lJMXltmuCqMP3H
PwQzjuuLMyGEnZBvCAa6uI6Al/zsOxCsyausuj4rgiQah9uWgj2kKzouUa3Rt7hnz9yqFBBoQ1KM
beazBE94/s/WZ7C+aWyVmkUoHDnWhQLeyQ1d+N6JWchT4vWHm+DRj9G697gZgroCllCPX78mMGhv
oi4m+OAHYJKkJ1G5HaqGYe2MwlddPzworQBTj1Bpsy97PAL145QacuqoO/b789cs+v/6TiVsqvHI
cJL/nykMLJN/9y75IBcXmR76a5h86r669j/X/aw1CsnKYVjzc9M9AQbwpnyplw4IVzgNouHhhh5F
Itn5VXQXM8Um2Y2JhiJjKKNBY7+R/v/G1kj4fnKeRQc75mq0CizUFgTL8SabzL44hNIC0u2qpSyv
TGLLFSsRznfmvRRKboCRiKjLJSiUeX+MOEJ0/E7cT6iejWsvnx73IwHLQkZnIZNg9jCdBkuW+Rcn
w3umSUnA7WKyW9SeDw/8qEHOo/c5fxyM74tmVCAguC6UMykogPBixe+GcEwuQdCEKPwQiG5MZX8i
t9Ry271X5igwIcARUCFXEn/QS70ctOE5XT7mD0Dcd+9hQj211k780dNEReIzrE6Ae1KHwHp5Q+Ib
LCQX8zkFeKQ7tmne04+UlhdrqRDU9WwvRIOlhYdUtiHtIMEUvrQ6hGTAom/QUZScRkfY9ob7FWSa
i8it3i+9lyNJ/xdQCfiIufViR93h45IUNx72mLlmoTjs6Q0cDh88NFv7qQbVQUnSMYrctzoPNCsM
3iy0eChMowcnvA8losC42SWHHIsHr/6lypm7IB98aDHoQzj5fqQ7vckCOzHO4x3RBjT+RuBzUBaf
fsdhD0V5KAfyfLMEO4tu6cSDfZxk+he48jw9AtEv24ltwdeSu5tpx8Pe1WWt3lZ5ncivC7LiZCQ2
l8JNIdOPZaEvSrlTGWHvTVTV4AtKjtMvP8/tOTFLEdjv9+o2M6QtNVTXgwScoHguH+adgsqOFzbc
ljipDUKPbk1tEeQWgTMV0MVETUKnAMKWfMqlAsDLFIg3bWujSYjnHJT9ILmPNOYw+w9zybQGyiUm
662VNXpMZYEbbFnguwGvmZ2OffuZjCCuJwURLXUopNqQlOm0fDs4xYhjOpDlcyYmstBzZHJg08fh
604evY5aKbEAcgAHzKV0evDa/WXz2uv1dGoOr0cw5PxjcLN8OUVVVOXiz3O/+YCl2iyP/4y86xkR
qKqCgwiohJitbJhrAFFSzgfdym2YFmRGSX1mtot6oiwkMW4kGfPkMPYBSD48q/uZEuj6HsG+URZx
CCi/lqTqRqh+J6OqPAFZ+EmoHIaL0M7um2JmsNJXa94SyxPnphpcksTSHa25VzQ1XNk/IWuX8igh
4ne+UdhWbU9sDB3F0o1Z/QLT/+I7TCLo1ui/X7vbetSD3ySFrKeSjxrHBNPOBBsC9DS7sQ2vAdZx
f2AJ7PlGf3T00sG6FlyrlYv52LHGJMzv3Z+BVnCg3M8sLDUMEMmTvXKNQrN+me6Lvkgl0I159Iam
wIgWIuR5kPRItwM969CvQxYxTmFwOh0i/nPuTbjv1LlVIg9Dpd5ayft1RpKKh9UR3mnqSTo8UT0N
6CEhZzc7vtgsdXP5BYUYGAptCfP7znhsLn9ZrQUNIdsp1wjjM+9d/FXjiUSFPrFsnfnM5L9U59m2
qS9s7/B8KKYF8fXvv7haGv4dkY1oOIol78A3aK2hxCmtGL3J+3WuNZviri6p9UXeh92JalFJz9o/
zc1zJyh8BWrxW+ScOI/sKEY9j6HM0C8yvf71cd3Pu/slXl5CK9KAgZulVIvbPHKgxXwzMYBX74x0
/jXFmwWTtyfD478mLHW3UUBHuFC0x1CSKQmdMQ7R9DFcokK4YzcUsUcEHmuIieyYo2W/0iMliAsJ
I5xvfSTtbUNkZ42T1LTocjalWmRBv7KkslZV4CrlyYufne3EDSbDLF3Rwc5MxchsE4nh3mOi3gvg
p6J315jstj142QpvS6kv4dIRAk94unU5n1Bw7hZWIOz2Fy4m/e5Y3NBOfjxKBvbuLdpqOZUIZp5k
lMHl7RZQLg7msmt8FPDDkjJayREA1o06KJxDCP70XoXNbej/idVkMmg4i+SH7FbAro9Cues7vPKO
R40dDi1gLpU1MaXxZVPUsKOZqe7pWyULZkdqrVQySpiBEmho7UcIGNSUGWphooW+k9F58nbvHMa4
EscQB67QdIYyUFBpfzp4Cwxcwj7bVxvhMALJviCOWjfe3DyoZCnhNsizpr4MdU9+Vhqn25l11iLV
06F9eIvNUhWeRmKr/7zG3GOvY4KUBXckeRz2dTuXZcagPsUbi1be4yR+J7ell7AOT2oayyqSkUXE
YFPoaNKEqW1lc2LGADhO6Ffhx2kGoBcZYtgwEBoGICYDbxhWm5NKag0oyoV0YPhCU7XDhibWf9Ub
oKywFauJrT2hDB5gQt3GggpwUc7Eyn0STmt21FkTth4LF40LOtfc/kmOXpmPkfKd+fVOG8bZaEZd
qWn2LVXJ/T90IneOrrEBIkAsLcjCgwdI3bODdy8CnxLhX3oeXrj1kK/jC4X9wlV4pKQBR7YGI8Hg
Z99l5UBxzOav9Eu97FCYAzBmvV4trfu715+Dp99kNYBa1ocfR6weJRFF1oZVpK011X53JaqtB8sv
FsbAolAimB4R38SuDjdSa1kfVAXwSPDZNdXMuKaHkFIPb4JethSRpaPtBHlm+r3dAtqMhbi2tnY8
qRvLSUaN2UxboPpf0dtJ+yZSHJ51LSXcb69Fan8nx865S5K47J5SD06O+9ryEkk4U85VCnKJlXAD
jZfGJ4uZw6ZurQqOrGnga479KLly+79BVFZRh2OPa4qtU43zylBRS5aUZf8gVYaPWYbfQpviDY4i
lmKU2/6D8HJqXxmpAyXwyEkHzhBHxaRkxGXDgs2cS924HbjfBy6aK+/ciz7/0rG48MNMQDth/Qx3
Bh+WWLZ3pCg/U58y7iNbbv0kHMXRBnLBe5HyRjqvHYFq+otiaSJc8PXnkKBLtAjEW/0qXP9Yly/u
c02F5Rc0ji6n81MKcZEnEP9K+zlxdzPN8CMJujw/jV2zlHZPhyhmebUaaNvahM1oqt9xPOOJwOG4
CModJRkq5Gz6ug2fXDjxeYcJ3725mADHl7h+0oDqcysNtzdEgLACblHVh7QQEqNs55Mtutn6aIet
PIcWyzwHmAnWILbdc9dZcbj2B7vqm3Eg/Q7wyylt05yo5Efkj8K0GWEZaGZMkvIQOIB4txyNi+By
FBtP/M0uhbHSjlPLTnLlZCGKwBSu5Qxqnu1Gmw0g1dhSEP5pXwdEQt0FI9I03dDegSuYCo//AuBi
sZ28yT7l1LKopv4tZJ3nNOBQgJdTvx446/2MweICWN31dj+B1WCfZ43Y2K9CFIq1SN6FVrRPqhib
3/npeQ9Tzp1UQfS1Q633Q+bshms6k9ERvcFK6eDgHFvlf+9KznurCRWJauYs4SpGb/HwIgYYwnkd
QDYYscjj3R/e0qxEW9VIW1ObwDdVerJMpXsVNgJ5OMc11oqWekaSP58E4GfbJz9fT65luOAlPZpS
ay5vphMSct0iUv+sfUtQM2TUy1L3mG4QM8LnTx8mxgMQZuahLmlUcDZb/NBDaATeSxZP60AH4oZw
H6z3Nmh8k6yrFeybGhExHilee1nPbHb4QgbMJeLmQ/7DsPYplarmTgUeHyUP0UlpS76kJkG6zpaV
SonyDLKrxajWg7dNbgpw3dxXmqE5k0XQXCPeohALbp9nanuVwSCP+3TZZeBnWiFVUwtwsB+y4sKm
GcyvzmJTu4C701zkY1fnm12qEVwSH93wGQiaTCi3eNgRqx3W1cG7vi0pgaYfTPjLXVoeKdppAMVF
7AbQgcX3ypxpd78tR1mPs7dAiMtccno4+Ai9ReME+84Loy2KMvGXpXm+dIXpJUq6J6JFnraqHoHT
MqgBGgjPcTgzHx/ALCK4+X53z2Lmlje/xZjSIfNEMx+x/E49MgFYSjP3VSgeMhd2NNSZ3MupEE28
0ga5fraQ797HC4FlV4vLw7ZxoL+FTWvatgxsfUKz1jrpAZF3r7I+sK0NqqCz8vG3iGZEo+tKpnEP
uUhaDfrVCSgm/7AdknMUSxC5djOLm2Mv82Av3Y2yXxT9el9BAZTxKGgVC3SYKPIFjS9z3r/VMZgP
0fLqrVfd6+38+YZvwe89pmrIVk/U88qWfWFr3MXuuV7XwT24fksHTWeCIV7RidJUG70/foKzQuwj
T3Pcaq7Ju4OM7/q0JHnqNMoC/QujNCTnuIyzAin6Rz8jeuKpfa3IXjrgGesmxa3Hu+AbVr11nX5/
vNnWjrvKcTd3T0BXVcyR2h+/hAEqtJH77RSyL9rnf44JSlEneYpb8XaSPOmGWmGpUJ+IdtcY/Mf8
7DeY6jJyO25ZVHcQpXMjOKruge8PuwQ2OZE/GJJbQ3pu3Yl0uc6hcQQVGDK654xPNzbFOOUH9Kpc
Q+Ez6/H29EKHuYrje5nJjCRFkDseB3t6us69xJnfvYhomUQgSg2n99PxVSIjLoJcqMBUxhYx8bcW
9inA57EP7ZgqVLCRoZ7K7RBE/gC6BPTiFAKQANf0wONys7DD2Qa1V40odZFdjGLv1XcKoj7KVuQl
dEv3aYZhJZPCwRmIs0Ek6M6Eh6LeuSpizR3d4qvpzgrvGHxSiMFXiWKbrL+sDZpLRxDNzDeXOUNU
Q/KjdYCDCbPbSJcnhYC3Vty86xu7Jxk/IehXnOWN0N1nOllnHhUQZb5UKabidBDxSYXPJAiNxAp3
sU8eT9yY1EChBNHYtK8xvBaoDRuATCs9rbiFyolXe1NuxIT1jbe0tooYcdfPxaWvfhiGr+26bY7x
0Z5n5dEde2+dJs8pnmWgfDkdCr95EWcg45q4FtVeDyUBnL879bD5T3Hq3cSCL3kfmEJjkHuTuoDF
kr64lMnBlI5fcyQZekhP15BjInKHxB7lPXBc/mYvTIkvKC65tQMui2LiSKUXuD4EKgiUkJD5ZPpk
Z6rAzF/PKf14dVqQEnJATWc8wgx+vAXQQsaivBL9pj7zkKRBTs5lztw1rp4ZVkTNN54c5XQI99P6
DZg1daY/hiU7p6EpobZW1STcYX9ld5zHQZfu4YkWkN2BXbl+PvsDSkV4B/QKOu/XheyxCimAgtTq
1eTwS7t6e5Q8TL5fNsIAWvEEvNwaFCr+vi9XBPXzf492aa7Ib0ittAyCDAR06/Cu54jPw/MfS2X3
plkgNrve//RSfqwAH9Kii7A2RmOK6/Yo+zP2Q/xTYhTn/ngI2cf13zBJsyuK+ROBtbykvg6v59zI
0FWp7qRVn6KJcjiZHbPAnR5rDUKFttU2tPpxZEUBI6A9qGzDcc8grRTR84mz4Pm8d/q7RCIpXhMY
p3x3wvfnKl5vu/Tc9FuC41rc1yd/Rl2BM8lb98HTRUHhhUrQCNPi4gVf8GyyLZw3Zybd6IGkGeg8
opOuvMhqeWLh7wlH/ExXv1UaH8Qi6H24UQ7+TbImF/WFo9C6i3m0E7ohtCVddjQbSPSrmXVb58Ct
ZJ4hiFBEoQyaJnb8XG5Bnsm4dUxgfZ+kxqSR9vsBQZE3XIhbg0yuFwbYjM5hjt4b22a9OkPsUJdl
23gkex7+V7y8S/x3S7JbumeSwI/tsP4TbCzvrdwD7caeGudA53o2wBiw2i0buSIhHWsyLDPafwm3
4AfogBIFqcPyfZw6gFk2RA2pAwTMPi0f/XdUL9MHd1qQOVSXQK0E5+yGPlBjVN/ES3XsBrbQBHql
NzwlwuurusKNuq4muqiB3JIBVkjVNbxLIL8UADI/Ti33znD/1A3x8y31Lk45szKS6oZhyTKVw0IW
C2k2XD5KLTla1F+5/96K+VlwLeD4PYsQYJIh8RH/tumgNTebYED+tBt3nzu5Ipd1iDTlkl9yy5B5
+rcY1nxWtSisJvt6bvlpE3j77YNSaTjdhVuFvrn4ZlPgG6vZele9oNnsoEy/raemlNoEkkhEuKxw
wLwT2DXS4yBtQywdNcqhRLyx/jL+Jwemar+5X2DxedC3WC7nw3DshsAWqMO3Ih0354ET8ooOqRrI
vPY28wYhN7DO6ma37CQ8BXp214D4zk1pXM3+AU+UjhD7OLt/plz/5R9Pave2B5WI3QiDyRLKBNvq
0RyGhbOgABZ0mgy6SKlp1zPuh8SixdVIVabK5+zY2OMxHdMx6PHJPQKp83Jd+tBP5ueDMQ6/NU8B
EJ+AEtS7faV6e+tZhEfmHSSpcs/F5FB3Sm1HUpfpmh0ElHFD4g7He65p006/+cmau1Z9DwnrSRLV
lseW3TkoWoouGzAraeQrXOZrGDkBpMlmhldR3WAbX1Ue40LI3j1nTH83apBMpqFFGq0AKsN179OM
KTLYTCO/sNAyYjPanWT5bSutvNELgltaeVJJeq3Cb9s//kMEKdxurD1xCU/syTLIx33UNUCOXwne
LdiTlRF5RgACqyl/KcUpM1vT9l4okAy2izttBzv1mudi3Ory/Q+FYS8VD6redf6q/8PKzPgDzPT4
c/FL31PcHrp0WmW0DLK/hgYjDTkxtb37RuZMcJXTcD22LbiMzi55XgMsCJQeqOWrOs8RofgRh0qp
mcCNVECasjxi4ODhTAAKwJnS6Z9gawP9H3dWu6gApCW4PE4WP7xF8AWD8JQz8XSp+GQy5RFhH1Mj
D7IrKgYv5uUdy5QDPUvl/sx+I2ggq99DB0DSxhtEX04PaTy4ZnQ7lhRclZjC5yqDFzeA7LQLCrCO
qO44zO+EqgcggMz5/B8aZZ788xw1TlH69Sz4AkDuPLGq6LiKWNgskAr58U8w/yLwEWo9BrFJAPXb
5PW5bzk4YZzzrFkIAuAjYUG0xA6h4K79urC/GGRqXPS+M18jbPIxLzzaBnDaxIkJI9bjwklHVidC
DVhfzt/fTV0gXSeb7VKSk93Datol197HDy74vZpeXeh4/vXd3kLD8JcAjojhdsMC/Y3gu0M/QX/p
j+y+uu6IFIR+wEktqUWsOoTNHhaSahoaIFGPPWwjy2dU3rijpn6j3T1jZcRyFKqpKuOwFLTIK1NL
LoG/qJspqhlZvhF30FzwuKDUYdWCn2diZPxkCYu+yFiyslgTowg2ozSIifbYQGPJukMhVEVASdFw
hCAdiqt+25xlpgyCIT3P51WWunoqt8V0PXt00ep7H9rOPP1FTyL/4/VF0nghNvI2e2Yp6mRR3lAl
ZPf/5HrFnGf17zpW7YDjmMKbcjaOePI0sjkzvTeuE/iH01eKD1ivDZZQcw0hpiHiOIkHIgLPA8t/
S1fgRMi8P/aTzsRi7vVjN7RGqj0gMELoUBPFRvxCZuA5GpykhyAvHMhQ1YF7Oq6/I8RTPQPBDjUC
pjNhD19TCIbibb+y0sHgogjpt+Xap3mGjUJYJEQKEcoWiRlV9j+oArZXOSr/zO4rknQBHdyTMd8u
vwImtuBG7tikr+M0VIAQmwWBIBShUQd2ZEIVYjG2hh7m2Zv8ceZR3XAOMS0Mj0r1M4ziWYEFk9EZ
MeusZ9viSZhm6x3nmf4A+KaBzVsLmOWyizNwJ9j4bamAac3N8DF+kd6IBKTufx1OoDhkg3dzieLt
7w78y1lT7iUEf6bZpd3QHV0kNvb0ZciWNFfhcDfBjirPPnegV45N6sojPPfzbcJBTpDLE06oSm8k
lYpE/UtScxAqnlZwVu9Rz9AF0EeAzzSvlhfzESoIP26EszmjTG7ezKeHgINKFi4OPuvxg1mcPXUu
eNYIzIO+kPPCkKZ6al9qMS25oCsXy9m4NMQ8hltTt276c+HPW3LdZaLuQpSsb9agQ8KcYxu+eLxX
w4fiW5BCZikwn0h9zOd1sF7V0jcG+sxCkklIp4cTWjbywWvd2J4i3EeqC17KNgKv5QmO9HIL48bz
kRPuUTYHasqFxPJjFMNVmzdiJ8VEg6j5eFADZJR5XT6lWLGTGMBtZ0WNRd6ChtSfs8Hh+kfPmcr4
ZwPdx2c5YffS4fNMalK7bhfJrj5drUXQBeWlVMiGKS82IvHottex2KRX4ctaE2BVbR9RHFeeG49F
YlAmn7bekSzipycDoop0A9cTj3h1TOzkPUXa+LpA7/NflitK0o7pe0Eg03IdXHtCdrOcPlWtktcS
RE8cz5ISd6euxEw3N8MUff1mS6o6Wt7eauERfClwvZYIdGjEkviAkAt+cDz5SjNmR9Qw6jap4zg+
A5cGcBBbhG5+NmWKfm4mGftj/ctLBN8ZXhf9PHUvJn5lOJ8wIaOJ93vFDSswswWTiEAHcR58k4CT
mGz7FnpZo16gaH0YhkG+2YTz+1PuldzZkrfwTYapkaZ8rcWUeLlPTawWvYoy5cLhKzkGPBvElED1
m5lhMGefgy3Cux0dFMLah8/YhtGrhK98HiVPxrS59nlWT1EbLAu6yyDljQuoa9H+OXCdgQGNXKQA
QxsUZYjWd99meREeH/+ZI/9GqqPI7ttYUk/SQ83VajreQVo/drs+Ru0z5osiDqwc1QMD9/mUmIsB
M07WyMzNPa9gcf4N/3Or5nJcyoSAU2Q7sQ+t/z8hiWPzYmb8fJluBe8I/CY2WxFy//Ouv6lBH0mx
8RA92ZLrqBQoq7fgntbCL99jZUWHwnEWbx4l1XsgfnXEEJ0K4sNj4vem9DK8gD2Gs1RF6nUe0lLV
Vl2CvragaVioqrYNmFBpQrM7P6Gto7kNTln8dCTPn2EfSO+WmGYnKAQpxBHSm0mh7L1QtHX5rlSv
xijvqm7RL9c7/vMk+bdbdHteoWjKk6XSE6jp0aUvlnf+YNPJS4pOJNX1/Nj3cBFDW7e6Nla+oxte
kSiPW4faD9YmgS8uu0YXE041ixo6OhfEQ4Ubfu/iEe1mfJ0GDSwwQmJIIAwWv2/XVDPkj9/uEstl
qeffpi3Z/f9RS9meGO4Ch3I9iIaqErMmI+JHLn0z8BGnOWvGPY3rUzPkZ0qWUWkc6XHLpuHq2nz1
xfuxTQ+CBE8+723Uws/k63MU4AJN9v47Gig2VJYqdgHD3GV9ctS1Qyy4xiC0A9ZkeZPg3eHbEG4w
7LLYeqFTWEP2rbZ3l549torE/oJNSCyBM++1AfaVLpKlZpRkbSprGWH9cIX697gc1Jyqezd6Eumu
gSwmGtzjOuqGGIYv3428RC7d1j/a2Ql3SiCeIQ6fqkq5XNddawzlJ6SVxWmoMHFmOMc/kHMKCOEr
rOZ4Nx47BMiIWLCdE4bMi1iy43ntFbUIhILn2I2aK/70uLXS15aSdr6XOxuwET3SmAvwfV0P1z6d
/n8qlfwCp4q/qjx8+qTbQowJaG/9as+TkQQ3jDqg69thAX8AfuLg5Nj80zAmwIm8oEW9NFKVY8vM
aGwBIEfZ74aZ6CPCEU/e9GKaSSMcbTZBu1TNXEaaAma0eHVfRhXm6rfPj9OdZxv6qrBZDSBLucpM
8LJSB0ZA55XktMUNfPU5fb6Z44GNZEPuy1ijhUVUKQzs4SUTDjL4R70dxbWfBTfwJ9dnqSEC8Fly
tVuDDD/IJtak3qXcg9rv7XHDTJvTjJYxxezxLJaBODSAuAYcPKolSS9ekNR5/C/yqw+3DM7v1b+s
CGNQ+n7+KUg/a9URxkB4GxiSCuUSssYMBQD/TyT0ntUCvTeFTTMtupOJbECpvAiQAVSpMLztc8qE
6tyn41rnVFPVH2j/iBlL04hyfq6x3H1kt696rOiHbuTvk3AAwiz5BaitqkQU62/igRHfD5BrWPJ6
BFzX90RlqbJQP/ifzPNwux1iGBKRWiI92J8JPLmIlImz/8zAd4Ic++HEx89yo49j51NUtdNnVlpV
HQW7ZLgZ3/b5pN1csw6oGA+3SWaYs/hTwAsJ/b3Fx/E03wXr1GEMGIFctiKK/VZ3p3jBnqEv8sqk
nLoJltWs2KUYYlOHJeuUQ2AjRkL7vKDw0zv6nRE0RBu14MsPdQG57TTvRWo0O6q24h383ViXplhG
stHfvTzdud3rBlIPNNahUephEb8+t13vPY/IX1rhJP4EMBsdOqQA31UIgaROHWX0Y3vJwZiwQPnr
KCxQKm6uhH8WEat3MkMsRvoLQ4nAMeTD/DJSUmAo+erb/UI6bUqrctZ9be5MnEi58NxMyjZtAZ/c
Ssu8MU4nKbGQIotST/z/UNuHciZ+ZaIvdhCo/ChU6KxDMD1GCKvW+BnWeB9pVPUH/TJE01uskDHr
GfLl+XOWulfaVnMbajm4djAONbXcma5mzqUVijzxse4J6AuL3p/klY9oGT0/zwWO+Ag+t/QDRpdG
wZLWtdSDyuWfvSie1XfvergF2M24BEgDRK1ZVNXarXuPk2kp7iPYJSWNCCwQTwu2LCcPPPWOTeTv
Kl8CVxqpEpVIViGQZTmf2KVbpPZ6f+4o0xCm/sM3+Yss5f/CLto5it6jWW53NMTem0fo7YK5X5Ig
XDjTPFSb0vqredMdG6w4NMBRbD3ziTlUQx4jNmRTX3UaO+kGZhs/FX7W2Xr5VZ2FpbtqsQsugZr/
JTen3zaktUHlfh7k1MtN7b4oZvbe1K2S/PK44KZxVcYGNQwIZ8mYrmKQG0pVlnstCZI9i6SJMr4F
5RgqvbY4U1BpOVJv5/BUB0yIhpGf4+QqeYOG+RrY6eTd5BksRC52mlAQ6B2yFn76PdkxWF3pk9Rz
7vXDWwJkHPti0/xOBedCmoQcK/4ruEz0VXeK+X4hBLcYq0Pu4NiT28yAII/MIE1+B6r3oSh4eC4X
jekVQA72OWUHciXhK7IW51/yiKwDS5K+bipckrDqVfJWml/c6l9CcvLBRd9CRCU2ae2xsh9hAxiJ
+pkOREu3x92NVlLO2wm9D/uHQu27TMCIZJ+4HVcFNQ58l0C5B9L2c95il/JPMpZpNic8djjIC8Bh
cL2ql3Ysv8oCBYsauR2hKc//9ZABxLLGZMRqVcbSOcPSGv0+eXTBhPJSbyHPGY2EySX87klx4NGp
lC/E6Lt0lqa0iYpUGAYRkILVZCOlfx3jLtXeObyZLSYnl06soYlUcYPxWirVRtT6UzZuXL9idVGE
8vXVUtTBJLD0mCyWOBRQ9/ZpvpfV7lbAAbHnHdGnFF/DeXUBj61Xp83cRtm6VnXy6ISCf2NLGll4
AIgDlshh1XMu+Hc7w1lk1gGghFCEu/wDz73BFauUZI2II3tT7GwIhDy7duuZbsMqdQ1DQu/DSdjm
1RF/QGLm9wDwaRhk2TkuKwv1ePGt+qgw1xuMTT76CroRguRZfZZhp9tszcSC6wimufFLsnpQXJDO
zm5RqzoMgOd2xyU7Kwgl60S4wyCrAJwgGB/MJtkbIBVFLdT+9sDxQzBvJw9eAf4qXH1MFjDGNKxl
ZQwMKq194+CIxYqb/eTzERPU+akFbIkKK5ZDqjVeRK/rP97OjPLPLSYGA2RX6iJlXPgd+KdJbICP
5hepgyuD1Xt7JZ85Cru21QLQmxnoF4+R0TEnj+LnZm3wgIJXCKuAWOrD7EhFE+oaQYfc2t9+Spq+
ljtLVaUam55x8fh9GVY4qEnvd6egcyv/sWEAVWZbb1RrltjpK7pTOkMJXa3rm2FcXDVu5DLaikdb
UvAIr59K++3lSlgOIF6htuAv4unwgIzv+Zl6z482Nr/0qUU/FH7V56Y5MFRMZuOxJfsRr69759Ty
w23Cp9Cwpl0kDk2T5FxVUgEYje8aho3H8k+1g1ucLCV1Od8CJcMxpkJoKxlzVWWmGVIC5pzDiX9v
z0Gxl1PjuxKSBPJkyB8agodmhrxkYT/LyDeEAy3Kk0e7ABkeM87tZvhsjdPRjRDHt/8no6lte0Q+
zESh7MtusXp0sGHXgRNrqZ2j2ngnpSoeZCgBP+J9T7dZcngoq1+LykAC0CVaMcqinl5RDAI5x5hv
X7Tbr4efj7ATrY9DmsZJ0TXGjSlKu4HkQ2kob5M0Aa39tJEMPfrIH9Aqlxk5zjufPRULn0icCQ88
Douw6w0voyOcra4crrHfQX1t4tbHjYbZX8U1QSBxEDzgBiN5BZVOzi+ceO8Fubr/L/v6ZQ1r2fHF
jPUUqKIn+hYyZAGd7VrDlMrxoZ9Xe8vzHgAGfBEyNW+27klL6gKhpMmoJBNAvR84QUlVjYSBdNjI
wOjynshPC1wD+BIAe/PyMScFALJWZbhCB/zrujb9DIg7Ewut2/gtMyF9Wu7GCe0/AAAXcBH1eldc
GdWiedhkgz81eHA8uNdlGkzwEKlUhOdfMEK2cIaHZ31Dn4NXwcEPo6CHTyP3AgfKSI15sFtBhltC
5yYOGwPyAVxccPesq/tVY3dXrY087lYA7l5pSn1urwySXjeBAdlBxgaLoghYLCpXxG3FMX06fxce
ljP2PZZYa+0P8o4bFtw5wVnRJnqYiWXAuy5nSN6XBbhseQvT11sPYuPIffL6lOhmP0tdTD9N9M4F
6MWm06DmExUanRblCCxhKEVW9uGL8BfnExCNnK5wleECuaTqq7cRs98Y3yv1MRZE5yHHDndrwBB1
aB4nJOK+YhNJYDY+fLgwUZS92b1HREEPemGh9ZHymR7258XOaa821M3ktfs4ymjIevBelttcPXQj
mmwXsWyaY+HOPlj4zI/nHrC05bBi9p5S3czIigFXYW2vUadXLJmyxk4rpvP7qCl256/8aEvDx0N2
i8WSopsvXW57k/pfRNnDvLI+yZegZIa9kbThnBQN6ZP8+BY/EHgfI4Ljq29ytOPZyPySi/hGcNtG
rNdwDVjWPmIdgXG8txW2OcXmAGdvuR4qyYlunTmOyP+I5tXeIbY9jwM1hYzrSdfPFDoVO53cMPoN
ykM6ON9rZKHT+y9Of2yvl10CUVxfW/dMC+jSU6TxSlPUs1jhLsUZP68IdF3b+HaN5DuU7mzfSyjc
9CjifRaN9PaiLptTtzEibKgwZG538gMPfDHTFDplAs60V0DeKalV9qfSeEVcXqWteiA49bOkRLP9
KoyGjRN9DQ5w8aQ1ku1VA+gjRNP+Su4NKGlXUveEJMcuTQH5ywOz1mp8oS11eqyZBn7kkZOGpOLC
VMb5dCxaQ83jF1YuGKEr+ra44d45yT4UWWZUaIC6V4TwmbRl33DkYCfja1pD250dFnJnaO5Flq/w
Yt4iiBMf2Ne0boF6WyHkfVxQUlOOMG3QVXOHX1RCwNp0C3dAnrFCxkqbS2J7lazSL0m6fLTl7YOA
LGbbZJknLWCZTCy2vk5dXANIa4inxFIpAFBRHjEsWT9rgsa5jTFHjP3MxyPhgGPlhdRvM1+nv2W/
gWsm9XppL/68l1z31/sYDZmAvfQNAZ/st1I/thZfDIa5T2CtPE+/pwPZXMlC5wJ/RGhQN4rUKjwH
L37gAsS8GC8M/t/wobM0wj2Ip+fdzMuUIBvzfxIFC2ooMHGHsMVIZmtBur2+ho12rNqSa0Q6hroO
mLyhGf/NSSzoGQ9R6JQ0IUFi+TCya5PZCfBdrdSkY0eZXEHyOPc/v4EalXR2kksk1+GApiM1b8Nv
oNVIxEsDWLXGaJng5BMKmVpJhryEKkeeu+YJKDj65QHxD+WELb16VcNv5EB2HvnRl/F8jt7nJYsJ
h0gexTFRX6dwp1l3bw1kUZJRV2eD0paMM7kTO/c/1KeIbOvbk+qz6kL+p6HpqQuwGRfn5bBRPN9i
4uxVdx6O7aF8zZ9b9XxxAGZUaJEd+B/MVZUyUUFzhgKp33vCd0hVCZahEgnuvRZD5ftIyHbDXn6O
3lAdwoP5aeNP/5eChF6RGA7Qj7HYFfUwSjtmuDyTiKbSLY5qEL4KhFQV7bidcaqPwJj2sxNQvSk9
M7EnlEXG5SMmrexZ5tr7XmeoJ2ZholHbsr6E/u+cQTLL7Z1eu6BEcVF1nrUwspeIL+ghyQ0QJYbw
YWr28KfVbj3946Hwvs2q91TLZlk4gQqLysauSdplpJTPtBH+8MmR3vLhNagk8gnnHHIfzFwowZkL
bQlXml4JyjI/9+/pbZzZrim2hF/R9LLPoGCbXJ4Pf58TNATzI/jOy+3hxzW8YESB4LtxKcphqFyM
nuYEUe3K5caDn9Hfs58Mav6Uk7xTvdZ3uG6E2a5I2FkTl/jy3+snnPxniMdcQFPCo8G/oNSCh1vH
HxIJuPQmds23tIKMqG2sIZBQE6qQyqRVjo1E3tLJpaLc6Lk2V4PS5bSkY3MevCoqv3GYNv4ZYBcR
Jrs1Ab3mYdTHhjqEDoPIJ/7L+Nbw452OmR7IAIzFNEh4LGAN51JISaYce8nmNLffK3qFSFhUuFh4
1SNbk0WIS1BQQA/cNYCXXQ8xto+foo/vMlb1JEBZqrLHXXKLFEoGjAKJh0Vp7UevWDpkZiOi/QCI
Pl4d4yAmpa3aJyczqTBKzh4OAax9vyPcrvsJ+IyeO0eRKA7ERMqQNUP55IFl3yNGNd02phOMCwxg
EjYRb//JkY+6k3wy+aJpFEauWR6ShzQ+Eg9UrjC+zKa3mgYXiz2Ezc9w3ve02FLcXdyL5dl+70Nn
KXZasx0w1Qtw2lo9US+n5svCvHdegNHsRjMxLnVLDKui/w7gSmiIrSCOXpPTYnxosayZj02UBDEv
yI2MP+n96OfUCxYzC05PGjCH93DCT7W4LHVKpJUW1/c99VvMNHCJy5yp6Esg2AU9NsdBX7YZ5Jub
NdlqbAYrqC4zyn0nlY7DyCAZGTMfA75QfEzruXiadAf+k9RXvwwqeNcl9z4BjdDQS5KsyylLe1zn
tBtMCvY65yHH/R7cBOGGScUsfFCnVWXbRHi6tiUiNYMeQnlXyO8h4lmi+SWAQ2h/1Rs84r23ZtBe
JcHaA3AJpK1gt6i2fDghOmIKjCf+rwgaEGwISCroChkdC/P/3delGZf2uSC8RdVFAkGbWw/1SgRs
c4YhEhzxq3MSR7KlETzWmHUIJOXBmfr9+Rf8WPmzYofH/0hIhxO8kOmIjcPqpkHMsVhHKoEzFHZq
rQuyVeuGt+Vl5TMMWDvCx0HCgWJa2NS0jYPihDngAFl1Ld/6AIRUE7NlOfFso6zD8IQA1XaHC+/f
LxUYR2B0uPqshj5gfxMAOXdChcNxVAiQzOcC0mNX26m2E4oXdx+9+O+JecCiyqT/GlmwOdr+XlKC
667h2m8sD1kO21Kg1bbV+wf8Czh4IYEEwfvz2aDtlIIOB/VUiUb0UHo2q3IWh1IEjbcvqsWpkEqO
fvzHQOsLgSNvx1Ip8JAXclFrd7vj4j9up/oJt9jDpy9bjCmW7z3w0bQl5xIGAkPMoUqNKDrExcpw
akcaSfSjxm0FA7TJZJZkBgQM017QZ84SXBM0tnrtUo4eZWBVl95KlIp9UQM+E12fC9ItFk8wrIpa
0R9XajkwEawwiWrU1NOd+uWr38+uKc6PN7rQsWuAKMWlI4UyVJ+40AUbZnAZci2K2Sm6vHLZ6spG
1v7zdYc6gfe/yF5fy6iFdWSSyt74yJ93Su3u/vND0SFWzm8yh8OaaB+ByFFQdy/p8QQ/LwLqYj4v
2GtyE3686ZVzLvt7a6YNLMdcNb0DC0fyKobAC+42aPTOOral+MDXVdAKmtzwJh7y09odMStZBCLr
33zRsu2C+BEhOROfHv7dHFxcerZ4/TcyUrtUBKQyx1cSeLAtLOvhqSGOl5KcAhQIjZnIStYB+5Yk
zXexYUZHY/syrhf3rxxDUOVUvurn5+CGcNUDnCIDRyG3XiiErGmQ+nI0WFh3j4xc9z6oRMjSG3lz
VNOKE5qbKR2sfRk8g81edAvQjSZUjQOhl/nLytRSEI6577ctKFlK2niB9m9BRq9K9H+05PL7hNe/
aJeZ9dajeR+1MPR4uMW+RWrDYsn350HivU3f8HCwwSKaD7iblXU8ueLAOOCA4339N0mDvmA3exwO
boSYxuti2Mr+vpzo8eeAOBDbronovEC1uYeLj3NQW7v94dr6jeAdkAzMGD6LTE+hvv5wduH5G9Oa
PYQo7GakGcmwiFaSTxOvx7qlYJOx9EX/TsqJby24JDmbTvQtnsyx9LVk5TzcIv3IODItY7PigSKL
nnCK/+JMPevMhiSa25rdpj2NoHay8CSAO2jsVI0mcdyXoofVJH94H9VIbqHNFCYwC5xLGpEIQM77
OPP7RVSQCdFJF5T2GobT2AjLKXoVrRgUV86cw7r0ps+cXumX3UcvDCpC7ah104eGUuXcTnafuN1h
/RyNye8siludQRiGfX8mZpK+/y8PwNnTBhcb9CyEzS4beUn0ObqqOaHBZ3Sf1Ao5U4pnxqLnQUeX
ipyzjTb/U11uF3wLO8CEitxbrwOk7MBbB7iR/6ZfhiV/s8IYwIZNc2k1DNKB4HyD8YmEu61T/9A4
UIV6KIjqShixHVQi1MMOEt8tkkhYvzaCbRJ9tckM615R/NPA45NMy7gq5E5UPyj5TEkxDMzlxyDh
sri0aHs45AzZ6s8DAeIRWVcVz6Wiw/Ehf6kkayfQZxfsTAuHPJeWW7dCch2V8jMkq7iShQ+aBJNV
VNBq3yv77L94QpkqUitiTqHAoB8Rsx8XEBZmlCGHJwTR8Pk56rhkxzqujgtV+lhrKIPsaNlaFYRm
YgChPb3qdlQVTYrsQZ9qaIF2VWUt0iTTiZGwTR+WNbcEpBje3zTBIp1HV5QUwx+yT8J5/IJZReZ1
rf+sPEFxCzKVOpqVJn/67K0me3RoNPJ2gadz8S1i9sbp5vaTZ0LEHHgQI0qdEE01cKcu8UfRGkSz
DtLugr7FOrQqKYrU1rc3loXYt3kKOCoqwyf/um87NggxlNX3o3E2cFr+mewZg+GJcIkPAr9LdmqW
g1MSqA5J3vWeoaXfZ4g/bR2b5CDvyftfb+hrlpdit5/X7nEQsZsa5Jd5D+rkpJeOpFbVW8rIdosq
vWjt8gfWsaSG7IjQTnMezNydeU5yfcpbFHabc92sg/o5lu6+ACzaR9IywN2DI77Nh/PP3UzsrCRR
VA1OZAgbGNjz+QfWwt4zLB4ZjkZAkqUFoJC2UyEw3ZKm41xHowFjWOZJoGnyIQkvLILp1rcsfy8V
/eLyon6QJVjRUDcOoiRuhJLgrqlXp/G76n3AXjNNBVhtnGhRpmQ0K6OEteQ3OBcLvH95C/fpF9th
NAclf4m7P0XBGoSXKacC6X5q18LfoGUc5CgH+4Lp5OaFcxM/0MWHOr9+PAO5Ciy+SQAW8BuzZXy3
FnCTwvGegk/PDsYA8hnQxOXL8jPrat2vzWWH5QJ14/3lBwWWA7Ujkp8bcpV7Z8sPK/+iDwp1h2/g
c3i9OJABiiPQVNA75d+qOVCONDZgrUbWuYgclMprgw5+cenxFbS8Qr2it/Lc18dpJhy7Pmu/Hsvm
HfXDQJjrF30yCLyW6v9LEYZ9FKsPn3XpGvSrNluIKOGfmeVsJNDFJyuKRwyGEcByENdjP83qvBGs
0zftbVPbfsGi5olfke0pSyTrJUiMdSa5HzIkRoqiBLb7K1hAVzxj0Q55+8MIi+1PFnAey4ty1Vyt
crWn4cG/UpWsy8j79v+AzvP/7ILI/wwsbdwbROqm5ll+ypNmDv68o5VS29tJYRD6WC12JMj6y5p6
UYdTW0mIinuzvWglOwvD91hPTWlnN7Pjrz5eo6p5ga1eQY042IjP8gSuTsNu1VxPBqzYIoi/0ZTI
ewVFDxRjmjK6OWOT69dVsm+nsa75vj+bwGej4fAUvW3m0Y5S0CjDQRmcNUT1GhiWQY0nHiW4m9Z1
8b6hafFDnIrf+aMY6Qco+J0M31wTjuflwzgkn40k8sijGZJXTlzD55mDLfo8srmlNYKKkECfncO7
O49Xf8WAueTCLx/B8B3Ezx2KB9lDXdWngPYGOcGHokjJk205ftnpY95J7den//nBkbty3yMz5HBQ
FWrm3w9Fe/oRSxlx6uTcu988oU2kIFdFH5M94NGB8qtU4p1fzOAm6Rbv+v2/8f/nieGmORwX8qag
95D/cPmQ1hgxNxB2GI2r9zs0XbpQ1AN4ylW0fDlUVNxOQc06gpNS6oc3gmsZWmxCuALSQavN65lz
nkG1lsovytCPY/BR4odGAioV7UUWjJEvpIJyAkd2rm3ScEWsWyQPHpgk7fBuDJCe7nSMMvXa6Gi+
A+icW4zGr0nPI4mm9aYwQbY+b14Vdd9f3NNnsj91cud/L+y17tmzI2mWB4j3szPf5c8xYxXYcvep
WuzL4Q6/XFmKBKbb5mOKXmIRfOSB5ApAuHUyaaIxAjhQwmbDNwmIC4keZhPRPYK7x66S+KTcKUOQ
8v/pmgJ6HPNvRu+qh+hvWTtr4QuOMbfwwHW6GnW6UwbiiUp/wYYZP2ztjIRX+AwnhMFukXmvfQyr
lHdZPVdnifcDyNQeh17LmejC7SnUZo4NxwESz9ZfROXozGvWBngEB8YM6F5AumikLXAMGpCMxf5N
6quQ3Ksxb1UepDJDQTrt5TsXnpCFb3gkvrcILlwjXsHy6StCqdJF8e/dQonZtycLYk4SlpVyG+dX
aKAm9zRoQtLrtX6/uqgUtdB0XOixxI9GGZ1y4l9jUGGBxRFtKZobf17iT5lgV4mQ40VDApSc217J
ZPPS9XBjb+rFGZokQ+jdPAX0KWek4qbTgelBmy+CfyrIVR7DSjKckjCc0yPTCqBiwJg8FurQVhlZ
ArT7zYnUGYoboClpGRRv5Y0DbaWXKeUB2YRB9Ha+PL3Xge+zaIDn/oNNf4hjF6cppQfN8u4MOGk3
F+jDFVR+CSehonuJK/PZ0AY9xSLpVc87r5nnwHTxOZJnHLVXUItnZKmvyhuNUACIJP3JEj2dz45y
LkUk7tVDM0L/5gNLB68SzElmHN2NqS3ac1Lpi174INOwOMYhnpapxpadvcQfdGYScORSfLj2P/og
xlxlxn2fGmOFKEqZjR8ioRsjU0IUGwNVFatiYrOtPmu41Xwg4F3O/Q+G/Hwi2wp0lrMJFtLC6aHL
76BGqRYWuHnvR+KmbDRaZtSqrvAXQ55sUZNt61hijdq+nInOEpOKIvdegRaVYhXkinMzY0OgXt3Z
fhaQOcXZguhYBWIMX4H0Gsb+uiRBPH1TrxkRpPHjiUP1WnZbv1iw54E9J+uFscrS12gOSMPJB+Gz
Rzi+gWMgYiWdv9WKUyTFYsJNmIJVXpbNV19ApY974BT0f71dKGAthzAenz9xMMGxIEyczaw4n78K
xV/so0xdU+I0x2LvfqtrjEInH4xsRStex+g3f3+OvbkBG5bbiT8Pugkt0KjcE6IrIU6nvh1wT8xQ
Zk6z3hOYPLqHYnGlFp0WPEm1T5cro3VUjOiPsUfF47MMuRhF03vckJ6si8S1kOYP9HfcfXFOPuS7
a2x8FnndnHU88DirgHEe/Xefa8jUbXbwNHYspqgxkcmjLLxAyvH0RBRHPfBgMWGlzxdX5bj8OkEt
Eb+SVnwJb4SwHNBB7JYxDp1kI7t/NbJIK7/3h9e4/epRZtuUwhJA36t7jFBVqiIGVPSKLLT6XDia
vjLxRRsSsHZewt/+VQPW6aV8iptNfSTZ56ijyeBGqev/r3tBljDIhXjeVTR6euVJYwl1CUSiYKGD
gI4UpJbfppN/AK22NcEqbNTgKYkiit7XG0XCgP70iZpNGs/1Cxy4j8h/pwPIJp1b1ThuyKLOhnh3
6dxN42io4bEzbHeCFVAoVCoNxl4oyC08Vb9KNREXkEsMhbShGBhys2/pODKF03a/wVw3XIRjesMC
PxfoxxqrtZ7YDMK9z49QSywhLXLluooum5+LuqVkmfRMm6Z57asKMA3PTWfdxMhlQ9Ljdx85847D
C1/r44wu6/lxIoY/ucmUDb0TMOeGku0mu/hhWFcAzsW8cJ+rK73qGfOz0FlmU+DMxwen+6KYgvSb
DuztIgv4l0OmGeua+GJNQ8L/ngyXLXXPx+WbtVb7miUdhvYr2oqR1Xn5UvaXZyNC9dg6YS3Y+ChH
/NwIKfbuCanCX4ThH79hGphxt2bf+2Z3ikqRhShiOcQvof+guyUnMjPB0+QDX0nhuW30vMTs75Pk
5f5F3j9derAS+U0qp/jPhmthK+53HNT9FNC8JpjrhdPjpiQbI6u9U9Q1Oatvm77g9NrTe8rJJKFZ
hdBvWg+BDPio0avupb5G3fQA0paSyoqVE7v7jDp/j6XvtCgMVsiionDlbjnl4ZAcFGLUXmKiNHbg
6T7vfrCy4eX/AYT/rpKDXKcbqzxhKa9qlp2lOD7XkIuyxaem8upJIs+hD97d+93wtc+l8Pe4ax19
28NjNjEi53SUBlBBoacVEF23Vnru4DoX216/UUrWO2bGLokKPRsPSIdY8BdKQfKUkrqFgrUK3vEH
kcAazxWNIVyAZZJ0Yfu1pFPrzBDy+d63rB4huCRHvG+jb++HsZEspHEZ8r+oTwuTkp8EiTbyVKUw
4sqPW+RjBdmG1ci+Noxa2eztwgUTsJ0eXdryBEKOvA1/0Qh96zDFAnNaS/dmJwkyt2NxRSvNGmLf
aetJJtoyGylH2r3e4+zyZXJwnEB0sHS/pnWfFTGKIhaXIH3YyflrrM/+BnkJM1DXpxIEHFag/jYF
bdH7/Ju1+aFxjc48RV8xSCEJ57FKocKhqauwPSYCfpT/rUWqVqq/4JWRphvAjaWPnHM4OGi6zqvg
swGDNXyLOy3wcisSjbuJCHk5GpsTWer/eXj74B6YMww8TfPul0P6Swma7kddFyjQ+RA9F/1C3Hfz
jYUIYk9ZNKPkfQpLlYjWuN8x1ARhxk1icnEKn7kcSlga3t3t2xbH4MFOwLfuCxuZfZ/SFit+zB27
7sQWOmWQ5EsX9MHZ5ahVYFagzPa4sAlxHj50T6uR5OPFdsu2cC09UuSQsrix/Fq5V9UGSVRtDeUL
6wxJpk5fiI0/hhNaYcubltR+TqiUq4+zrDC3ZTUu/WplKYGIlVPEFV79BXfTp046U3PuBYAHGJhU
luTAVjAQUMT2pUxF6zljYgSN93IH9G5KGkAuQ4ePfr0dJGLUpdYXRZC8CN7uVGQXfTDqm5SxwTia
fNnn/Wfbom1NbQQ669az7YBMwPtTSOKJR1MC7NuLJrLajpBUmP9TIfMFsVaGlpKFJ4b3wCzkoVWH
5cxNq44PBWwXIyv79MJfqNgv/+PorY7+WCDD9Dkx3P5V/dXp0MLyYLsOLp8kZB4kFla2qlU1Rls2
NggBR2fqWXTaSi1sPvRpuc9H/pJFDlUdJ46zKdKKrMYZqBVJzf32lWuOTxCx3pYhVIe2YpThbPVh
yj00Z78K8HUyBa/g3svzmd6FdzbuJKNly3JnNYFiLdV8IzF11NlKKbsCbxZpE98L4iomxKJigSax
g46fonVh8w3dUGRH8YpAw0H1tALyT3lZrsglKwW25mzOmBbIBbyg0uvlPc5CF4LRFkLDCKDq1bWc
qjuMWLEmfENQlBqnPuuKVfIuNdD7qKunlJggoV2FUf/eWZbQusWDO6KqcOpN1puDatBCZeCd/0V8
ZOOqueZpTZe0VIqIBeRjarPe96D67r0Sm1Xy2tO3L8gIc04EogRBlCZH3utw1dAhuBNgaFrSvW78
ndhFigQwA+13STi14p4jbCfbI0kZVZmayxiEn2iMyXDlq/mxcWNByL7qZbrtNHUW/9iINUV/zq4Z
sUZthop2OJYw/fqsbn6ShbzOawoMc1JvmWf8r1VW3NrhDo41LMBMZ8azB3v2EflL++12hZf8eSca
d/6aWJoT9FiUCS/dW9FpF+rwdiul8wdQBLHghsJ2JFmbwytMhmzSUtspGHKUgc24WD8ElOOSZLlc
qGoknM9ZzE3pycPyn68a3eHMTFyAqxiG1UkamZ/i2yG4FspglNe7yH5HYQ77VKFRJorARUmZCAZz
pPNnF7Yk0VH2nTLxNDm5BQ10gCl162WLunAVzluRbjh/5/e0eKssETzDxrLl1Zco5TwCvVT9W6eO
5GTfwqbfeEgBRlgiXU1m5kh38DwJrrfclMjLtqzpHYwZojOY0g6OY3G85Nfv96x8oG04f5mOJg6c
CWp9FE5KBUnSZ7B+ppc6P2JTFM9/xQjkk4gC1IOagzBHVy3SQakr++2SURS1SaTuznFhQ9YODlGF
lH/EWBM881iACXCWuvV3HwjVVgFFsOXN8MJYVWanTQTAq2D1ohNOqdmMTURyNnotLq6IHt2ZhnOD
WL74NMz1E6M8uObl2lRWT28w7wnX3effof4yV/+gwbioXIov9uJEtpRARwPr4Zro1uU+qG/LlM7K
R4xTVa45VrvYLVKT3Kr+Aksj9e+aB1DsI4cKgXAFfsSBKzuSsWe4WxVSzrr0wC4Npo4N2CpwhzFO
JA79w1dsIgf2P/rIqW8KiPxwsa+mEZU7nr8K4bDdjdCAS9H6NKOShtMT5vMNeLBliDhj4k5vb0xY
Ly73RhaOGv7R0+IEi/u5NerPlY9XLo90B1BoWbLfSis8kUAokC7Q9dyN0xjTalKcDLWEqoQ0zYEa
I23UpMr9O4Hs2D3+TZDnbeyXz/2PHs5FUT+naplQftSZoXJ5N5eP8ykvczQUbT1KTnmI75BQRAoY
UMBCCU3qp++tt91E4mX/VyjuKRTezockdCJrDwNndiJe0y5/FSO0fnAAO0dhFzXDPeKaPHT3se10
VkoUAOAdV7eOrs4Gsi8flZRhyglNaDDlgLtLtGLwyaxF6tylAvIZlGqclSMXEOXV9umK2HujnMii
tezpUZCujNid4b4jQwofgAhW4X+rd1Ke0ZFnvM3mhCJ5zVZxVCcjDgHmd3WYe0kPYklkMRzIjFQR
s5ajXZu2wNykznXvOUSgtT2CmePV57L7y+45kdBcJBJ4XIoDRO61OAmg47RIWmMNWUhncuo9awWY
LOlJne2qXQxXnYLW8cNoeQWiA9muZZhfoCMTW6LCGu4ZJwDBqocspAEp2sjY3pu8axBA1ZVucDcM
yroHehHAjlsUQoLCO+ngXasbsJC7+C5mxcqEp5SmJlW91DD/kNVTqjfz1avwqvPZTKhPniWxyqzI
YDKJPZP9nMlnnQjRmFbTgUm8FugUvCpq4UNyKj6lcinmfZrKsehGdtKga7YT1jFYk1Lr99thZHXA
tBbwnhoRC9HGCY8lSKGMaK8Z9xGv5ccbGSPwO/sA1LltKFrcl4pKfW1zP3ijep/Anhlio59ffEqO
Bye1seQ8ZbtVIT2iJ3fpSHYaXqt21gKiKdaYZAtPWUTfQYf9Zmf2LOXKPFSIyqr5j3z7K2PavVfQ
y3Vbgun6fzi6TYjJEYyIDC6pNPwzMpJsxIBrMpOfb2pf1WFfE0MxcvCUB6DRMuyofiegx0aQN1o4
6uXod/eq8cDgwbvvkS84OBl/sVBD4/Bccge4uMaFbvR1M8t6q0+NuzzxvpBIfXMR02Hn3CUq6ZiF
EnBr7f5nqK+rvwfDMJqvogr+5QmbPwhVc+nMV0M7vB/b0K2WPCZCv9sNCFJo8mNw/bDRWdem5SIJ
Oai8ANK1YmQ8V76qVWEeUyOnh/Uk79M/TCGKDC63TWy+Qs08x5kyAO21hqghlslhWGxnb3OO71Y7
Deej+7t0ghHrjljYE4alS6z1moArtPcuiH0RlVNdF4+qKzRY+B4x+sM875ZyEnwGbE6yH/aU92Rh
+sh5DOtnIAYuwuoHpbjJHiEfZA9xP48q667df7VvC4Jd9O8W/Y+39iwMALxu5O3Je/lKdddAzJhY
Pnbt88i5DyJ7xLU2r8/h+paLwLg/7Ht776SoCQ5u2xHZyuPPlB9jyLhz8j72jMoKyEvBLa7X16qx
rA1WcycNk2ZQCCQSaMxB5ckm68yzQKEEtxVhoCoavRyhHU9LH+tb2IMWvWvMuILeUhivfatPKX49
rtRzu957CFPnsTxvEVdezKrXtQs5rtiYP4giI5oqUfikWF7/9d4BcZktsgZGpx5UdjLLW+MIhwKQ
9EvBcNvG+MiU9Yt6WEm4SGOUfzYBU1ddVa7N4xa97ryfnudsl7hJfYZ0wrvJMuiKMmbk9Tb3Ha2x
4bBPVkbgtcECQYKBmmuTrqht8Z4ubwXOsznopi4GriPhBGboa8N3Ze/aCgUUIjA5gfz8lFwZ0Ogc
mcs9TIN9clNh0yWonwRd5MXJC4e1axD8fz9yRCAxJ+gm6e94OFcr+M6QoZ10E1kwhevUnTipKCRB
AS6QcGPLbxsaYNgt2l0FcjFHuKo1HQTrpqXl8ceSYIuV1xyPU4obanZIj7axkO/lCht4axJBXbjI
kvqj0jIKf6gKIx8qCbnjz5ehNcZBC6G3demkt5d7/S7D425fCw7l+OnYpcj1BhJaSFaC04NajBiy
MQPfjpyG7Dimp5Qs5hM2Mosxj513qMkpzr2qC2tymz3gi9KNuXtvDAfZ2oLDkoqSsmX26xNHQzyF
TNhV+y4N0l84KZg3p5tZeKCTCtKDJPs6woUyp9JadKxBZmvhkFS3flE9JIjF+R8bIXT+2vHDcIBo
gFmKLLJNPQ5TEAdq7xgo8RgQBgkmHe7msfY2P/7qbKdrP3MU+N6JSitbYl4bCw7v7ehVcPEzDyrh
dG1JtzpWwL5UvYQ0Ob7aVzFK3LjDlH5ExyuqZrcP1131KmdrzVYM+zQ30ITcn3e75kRBqI9wSH8u
o9+H1jlB7If+0z+kOdZF7J1d1znvMDY0JmT5Gl2hUwULvWxygoMd+JbbcO9CRYNgyCjNrZpyjUtZ
pbdP1rvecImcOTYVaUk5EZNy+GJ58I8GHd7SeMBfTWn1u/Q7TDZFFYgfZCcH+/Sz20WGDaJzRDJt
eRK7bqalzyQToA4+ctBtudJoN6QB6nDnTICfyqX6/bacVFUjA3rFpVnTTinJMVo6IrLFUaHZQfdj
KkwTqdUo+XDBefICzcjxlJTeGjmqLzO2wo3/o4BdPq1wIhnqrkaF6bRiJ4KOR7qqHzsXWn9lH6CV
8JSB20VF5VsgDAabkI/eWHhv4/1IoYuoXoQ28D1Cf2M1RTuOb4XStaZg5+EN0vzjP00qYdxYYOO1
vJXqn8HNN4Pce9eVygNeQuNIHsJHKMr+7UW4reCKXmLRG4Idc5fDRCgCqF/MWQhH6J1u47nu/hm7
auCofKoRudF/t9Ls1cfHOBZyTBZUMiphUW+iJIVvCUbDzvOxW3xxrvEMsDMewl6FrAY1UydyH0iC
f31HXkDV5oJhmc5MztRq86WVI1f4JxbbTXYBVENcQLmegbj0lrYJEMI4rJQrhSHHnWiefbADN4O6
om+4GiReX/398TOJJI/wQwAqLGOBr9eUBQfPLlcCfDsjSlXxaf2UphHaUUqlD3q7pGq/+An2cSP0
WU3lSTUyYO4SBq/7IV+SKY7w/K8t00OhOVRtz5AWwu5TyfGYaEzhoNBMaUc/piTuRzn2Iu1nOM7f
1GlFkPAO3jbbdJUBcmo6JdzBL0kpFFRleZYTpkyOTn1LX8xFMa7nYfmUFwjDTHo83UJ5FAe4otye
d6YLEL+IvLqcQFTQYA2KaMPHGKFnVOWy1QxXDXWG//l7YqzUX6pA3mBtPhDq4NhQtcgciLUHUpDK
1cNG4zqA8RK5Av7bv45b38IcwN09hUbYVNPp7LAa5LOgGcVJtlefKsKRBKC0+mbR5pAynelNHrQo
6CA2nrBOS9L3AIotMrTk7j9hjF+nGNGAZ6L1Lz76DVqT5Fy0kOB03YZugVnRD0iqeKWp4Eg6C6WX
eVidf/H7mL5zwf/L1ZGCw652+VT3sFgC1ghZ43zXbhhDSUTschyXyR6/QRcfKglBfvSkPcmEQW5h
elVAOOeT+oznDKqvpico5OPkrbdT05zM71gug7knFUjFtTLWzOVAmFg7TAO3CgbKkC7krZxsgz5A
xEAYW39v7efty9baV9dR8/xhOjXuMQp38pGiZ3HDKWu4s6gIQGDyMIphDazbwEeCT1gO8rf6uSkr
bbxqQoZL48I+GJcWi6/zQu2f6xrDIICVWPsCcW9kpe3qWCKEFPdkPJfxRVj4KCeMHYhUYeftxlMU
mRcQOFhQWdSwHYLKEX6f50ktCUJ9BCDl0Q8KVQ+s7daTYJkJ8dz70ZIJDCbL9MHvwXn/1CaI/OjP
jV/Nt2f0aSEyK/Ej4mGyUkL66wZQbSKJKV8+Ql8AhtkinJ4hFtO+PvgIizkzlkEoL0gcbt4UBXes
yRoRievUbOIEJoGZ8GaN6k1FWAnbFEwtfSAr3om0Q0uWUNhIfhXbsw9sRIxGWp0lmL9d3TBKhJwp
kTZGAVpQ/1KjFuOuOVGlPayO2XS3iHT6ag+Ue5o2gqsjZOSUoEMi3Re7qtPX1uoHqtotkFKmETsD
x+eniuOkYnEQBMNCBGXiaeSeuxJ6oTE9aUWXrxF5XG+pRRcr5RTX3JTJTrIvtLQ+NP33UwkSnF+T
j3Py5lx6L17N5G3I3H3QF60yCDHt27VgFbaRkx7/DZcVBs7hCSFLMoMKXKa7ECx473fd23nWclwT
js/2ut3TLB2O8ycvcdbsfpVwmVJI8HczBeEdOtewM8gYAJMnWjoW4KYVCstDF8B4rddS64/YcZL6
2k8QVWhvUa9Vod9kfzZKlSBJFCxS/tp7WtqIkQEca++iFQbPKua5TbKazm8xhqZWmqGoXl6mVDIA
9ni14FY9EQS/xS0lVRHJL9x9eZiHqd1yNDDTBrpqg1bLiJ9V2wurMM2AU7RcZjWIxCygI7NxCDTx
MSQJInw9abUzrTqBN3EjvOTSkDMEpAjGKaczYRD2QwoyQiS4SRoPj6evnwu6Fks6StxnbLCLmn5t
2zJbGBILcvFupEd8Z+nNl7UkAI/gXM6VoUk2p/9y/l0DjkK3yjc09e4n8vuKBKHYOlvKJ9rOa1IO
E6Q884OgYtgrWDtm5/Y8Oe5dw5sKmGNqMdBkytu2jpErR5Kqqw2rT3+XQ1dAk3f01H2dmHojYIGC
9jGSiCxljb8gCmBmJfZyr/U3NqvvUMQtVv7pdDLB8ZYE4okXknowGohoElbZZ5FHtrcnll4V75z1
rJ7KkHcmrG90pCokXTLaK0B3xj3BUbNFNgY5q2RtDCY+C8cIbckWWqVqghFnSWlGkFtb5n5GqnQ8
9FtLjIZFKrB8HwSvIwi/eFp0dGvbQpYDgyd3/qeM7/CCC4Suhxz8MQeM339NscQcEmda9ZBubiMC
D8KvPP7oW4dfPwjjcuzQA9Ckw2wZXWBb6eO8mZUR7l1XZ47vdFCb7c7Jmhtxle6vbNtQTLb6xFOV
KMs9Rb+0dKy+XYV66zkq2wEYSSwrQCxMijxReZdtyDKxobvBhOEjhs9HOL3s2b2slpp4CbscK75X
ELpDsalitMykapFJMf5ZeXH6Okin0wsBZH3WBfYkINxQgaHpl5Mxu5L5002c7uZoGaMeriKkOZqe
Lqfc5pILcPQ4CIi8vjErjhFutgxrJP63NWfQhGcZWCN/CXTlBL+IAx40JvNJngT4LaH/5ms25rmB
YGHVfKlpMuLFUiI+64u2uhDPm6NOTy0uat+CjNJURya86S/9HWjapSUZZMDUhuqleEtt8u+NXnqD
WjUZTZp2THKFwz2Cc/5xew8JB0MOq+ri1J9VuffWhrmP3nnEdopgAx098TuP8r7kf43tSgTUSUuX
177M159ptLnEhovjPM4dHaaRHLH4AfCuqMDzj+iI2z/PvB1D+easXPv2k934/QVW7P2yFhFXiyK4
exYNrKJZEjylNQzpZzkQbIEK15vB12Fjjin1J3z2xo/HoWlpJTnmtlgCfgK/nX2YzhPP0dSm7T5t
5bOSyZFP9BiNBkxxoRudNZyVr6hN0km/WW6Q2UnBo/Z0CaLHc2kBxhrlV70LpgluzlDNxhd+NGNI
kkj/100w3jgSFyz+8c77/6kg9+SN0Cb+HVKPJDZgPmdBKUZOj053ylg+JwHsN2T/Z5AcUS1ENuEQ
NESGC1LpMU0l5aBkdPHwYNYjj9wx/WmR2CI1rxcSCZdnEyurwbB9UgunhvCnoOjukkSWFF/Uxre7
5ghdUlJ15jVvvpk+OLoMMPKWwzFtSUgLLVrfUgqVSQ6RxiH6M/ljrLBdKa4q9ZDqO4wz5v1TnzKG
jOINQsf5otMYlKHw1+b2F+5uh4ltL2GeQVk3/2FnnBg4cb13vPwUPV4+F/qHYb4/GXBqvJz0xP5P
Kmkw7KfBE/B+GpxuSQ4GOvf2jKI3H51kOUHLmb/FpEy6C10ww5P+XQB2ufSMIMM8skJ/ENOfFbMl
2o9c31xrZ27jaoNRcAZqcjNyOKYbFTU1dV1YMGKtTRiSBroanxSyGsw1jAtXfJfza1c13kRIQIsW
eHwXEuPQ0KX8ACuqbWNpx6MkSX2AEr+9c3SNh8tLOE54UPval2WrshnHBd12Z9Ku+EwHA/kTjvVd
VG5tL4Jspyp8PmK8hL/iRMo2xPzptS7BWvSYFqbMF5QykYND2ZQ074QzjcPdWETCFjmh22xo2iF3
hl/ANYXdBiWWHoX/4c9eKkBpHid++L+ozMCoy8LhfNO2Bgd/eiIcEnlHQbm+q+lQf1WyMAz7gGE8
gQkcWLuIVkZYAbraXz9dQXhabqr5fD5hkd4T/Xbf4GNkqt6aw/3Ziu/DKYRSz9edMhVlbCyzoYaF
Ue5XYAUI9PrFwXI/v1XTEOIvdXNoJyELcbygJhNMuv96biPIts3ids7iMvfKOQ8BlvppQAmLLLEt
OZigxOnG/jFLTzy8jel1HWcvgSUzGn/vORIDsjj8tR9PNXZt7S61bR0vIfKAJjZY+iGLOlOJZmeC
ZxOz07xy18I7eQkMqaJb1GqV4csyLKwOcQ0dfpqUCghr8Khs3cpmH9yn4wIIlAHwOSuzwcnuyo7F
5inhFx/IGxmo0vftHLeOhYHT90EENyQFInzj4tZMnB44j7Sx9H+aj7gySu8f6x9sPNwWXZk65A0C
KPquPCIcjH68fZX3KVLqbE6zhOjLveIPo62KLxmzI37bRvaez05WNQbMRhwTPGy6ssW7Kd8Z0JPG
AmMACbrZomvkzQfDre1x0+2WzC7ibASwz++4EVnlesJrR/xcpkvHweHzCFJDCRDj0OWD2ZfPcGZE
4K58gBUMRM5dfdTLsZSmQand1Cf9Hs3Xd781Z28HQGApIFKDJYhgihULUdXdGtv3X9n5dCTGFySd
qSPZ9yU32ctatQ9FocW7Y/qxK8aIAWmHvAlrAuCKV8HTm+R05lHppcWNshrqd9KTXLCmQ4tZxQac
zob4+bGP+crNYKBaXV9mmyvldG/GfkhrXNzpKYCOoM8KuavbErDypCbiDz8bT7HffrfGPGwV0BZF
PROCm1ZadA3gWONuYstuEswkIk8gbEp2E6t1+rmtKiZ1ryum6Tj35Wdd3UkoXZpG5FJ/7qF/ISRK
u7IF4K/1pegNxvjLr3mSPXobuL0QmbUFQ++eFzcgD9lgOc0n1cIfRhlqUSmcWjbekg9DyQurJ4ak
9HI5RfeWB2jLWC2u+lslMpszVtrCm8tY1NfiuNmBp9jIekAMFRzB4wDAwhxRXk5vp6c3aZo0oSax
ySA+UUGlJ+cTtO2orYdPntt2uszpW9xebjSmtr7llanelhz/x5yIRBbO6MPuLDm6UFbHvftf7ZiJ
dZl2pSknVTaVVQ3FjwFO3CdNrVD+x2hKnSbt8RePG9VF7pMKxImRB1+he0jV9yRfhG17KptZ6yIw
2B+w6CQ/gYdxzfPbAVwdDJnsLB3AlVaZwaMfomjwjp4Xdjah26KArctgMRjqLypiT7nCVm7Qpvpx
gpeVst5m+4iVT6lE7YyuxfREaC9OfYfHJfk6442adW1Q59XQw6RgTMKJQwPHRqEVB+nKj5Fd8LO9
9a6otIT3G1UsXIBbQpgtlIBKn1icJIflyhvRa5fUkMfYYVBbomPqeIgijhr/pvSQxb+pmcFE24FZ
2ZJ5cHN6sKAheuV4wh3tYeLNaausnCdaV4GA1LOHynJ/JOmjuqLLe3Tld7eZLa1XEvtj8Kw8Ry6i
OiqYIWh/uLMXlNZzdBzIH656hZtfP0q+mUWIGTsIf42oMQK0Wpgk+GJrY1n3sM55+UtpqgEPk5r+
qBl+lmEkJnFUA3At9LwTKLipA5CzWJw00GvNxsem6vvfZtS9JahvO/xzxtcyLCw0i3frYIcoAy1p
8POerTLWdJRht/SUfwGhKWZuiNwvSKt5ZAQw4RERDgCFzoR6vrwhi/mbDNeoPcR58DTKSIPPeiTn
czuN0HJDIASu2MVtHoMj4CVr5rKMbgk+eJ59j40ailxRw75KRtEwmbr5NcUYmzvkxNKrpKo5kHTu
yZz+ryrcaAI881fbFPF3Q+zjzfjXxkZt7OKOTv6sA0dXTcekB+9t5fjwTj1hnCJZG6MIZ4f0p3nw
z1L5VHf0NZ70X1luCbamFLc6S5m7PHkWvFgnjZNFfPZio9mncqG1AeTnI6oBZMJyCPtvvohWGhTj
wfD85tgaGvRUadScUMEuAS51r0Y2FBHEmUIYRF9HTJq54xo3PcQQGGc/ugz9VJxNxg+EGXe5QxKU
CSJvBPbCVqXAP99sI/CkPJw2LNtQ8UlBopi9HePDhUKtD25J+2xG9ekqq5ZAs72NfZmCLcDdk12Y
8e8EOZgzwaq5DqBzFzRe8MpSzfJaWkVXpF1KqZJlqZaG7J2jjpU/HR8chnfJbZPnsdhfXv1MFBA/
02psRPdO2V2ouRpzHSbjH1DW5W5Anibth2gOAAuhgpd4fBcXJnYcWYBO0+QnhJXz1/IR4/tzU+Bg
y9JtwawCX5wEwcNzQJfJfi+djKLZuBkyXifJHHxNngkbrGUzCIPklvNa46a5G9rxkRUx57TVvg/W
2LQPUZNMpiWfXAqyOde2UfUFNMWKk6ZFRC8r9zRWPGL3l9HwE01SoSGTTmE9upJkDItkgCYpNhPt
c0a5zPnHNCQkss9FEt9n5GQTXh5tClPZZqh5oDLlcciGW09e98AJw5Up1mK8es0Xt8RxQknDyjkj
Y/9Nn+PPOe4iSsNrGdFnfVTFiBsmEDLTJs1ldF68jbQ5CWxxsSq9+iOkh5JN7ogaBpk16QsnjpT4
0E5qoo5YixjxnSDvyiFpY3Cap3q/TsvaP2GiZLMnNcmeNlRbSO7G8d7Ex4TFJBeRhSHYCtUdaF8V
gbZZnFQwfoswf3fsuGGhsTfxaFLlvgvu+AdxxBB0JZouwsfkx+oRiSr0IHzIKKpPfWW012okGi36
IYIia5oXqArb9wbKz7QzVQF3zC/M5ZGzujds40uvbov8F3NyY7Xhr1dWR0ec7fhAdYd4jNDq7cqa
JLaaQdmroWSTCKZvfNaa7C7a6K+aGY+EY7oxqg0KqCPzmyJQ4XVdoUjTg9OwmmP3fmdbRMnLkCsy
qZ+TkEKKzTQIDe22iZ18x7IrlDEAbWQ0TxklPpXo0Pfn8e4wPTGbEgK4BL4z6tzCG9AHR1byIDGa
LK9pi4SypQY5hUFEDfFKtEySfTZd8uK81pV5PuxDLeUY4jYRFkyENmky5FHEGtzaB6Gwm7egbBZf
dmksYT6cF74uvb8UqnVQnsIMzuRwBgbr4c/pQKV/QKTeGegUH01UIkE2J4qA+9f3cuQ1U7m9Iyqa
wPGGUd/WD8YNnbS7/L+ExtwdK+5g+p1aWke3AnGfoBjW7Z2uxnSzBxB4RJQxzCzCrB1RtbpTLPfA
QxyCMkloBXmMtwb/Rp/0htoSZp7ZsEqTG6Tt45eNkJdJbs70E7tncJjW6Rsn0W7XgQ4nU3TDMrPf
dvm1yeUSRFVsbRSfzUrgMN41C+SmGXcDIyAYzctL161WUPUyD+riwUKRMtRpQk2gFvPOC823GTsn
3dtUcbqDX8xjYV4UCBAm7wKYcL5N//OLZKczcoecLLhWQPwZnaRxoDZjBegtFgC4LobVYg+YiUJJ
pDNsp0C0apzhKEye6xM3Xn7LgJg79eEJ6fUxeJxtw+68QqoVeTo2t14xubVk+KmBntsF5dZHvhCu
QtxGRzpjfT2IHmCeF/h3EKonVHCO39WnAua6jVhpqrBtQGi2hMjbFKOqY46Me/ldU1mHxE6yuU1S
whu6HLCrdZMtuptaJjEpWToHkCo2l5WIBELhCA1YUPBO3YEuiK60lVa/v2627lFOQfz3edbJQYJ2
1MJU/psTjlisSI02ozdukVo/GYirrP2E3b0PXVmm4ROdTFt9IYBI1ccwEYoGHbp5YOe9OpDz+ImU
dKg/IGTspl3IGiIiDRYHdDf/Gc4DX0ccYJPynPp7kBC+y+Zp8LYl5mewhhuJONYyk7eOZiPtdJcl
FOjaMzZPoyTQtiAbnfPcDonaTu5ZS8J8eCgQRvuKM73vLTmLPEIjYfo3P83TTV8dTUIYDNpY1DBH
d95UeBqdCQ1UZIJGByodmG65elFgTq1FxaDjNN9GHGak6EAGKhrQIAbVc7+/vCUKQtJJ2b6U/x/C
T3OM6AQ1ri5uDQpxojlyzT5zpRxd/7cxbUuVgsHddhaQ26w31u86lK9AWs07mkg2Hwi092pRSaTk
QV0YIcanfeKhtGWXzrMep7wtoqv3OatHtDzFW3+NYKYxd7fR5Glf1/t+gNSQiTGKxVByJM1zpHXK
AoB2Rj9KgYFn3xxxZW/lqG3peRdZMYxXDDempT2vovn0wM7FWDVyxbS87v2GeXnoANMx0kDVl4kt
aT2Gjtt7ztnPEUWfTVy+4JOgXj3yRvSRqIVV0we9eAP0YC8KwqT/zADwxfke9PncL6cVGfk1BKyh
3VaFiyzNvfiTWz87tImEojMhNI++nOU5KlqV7joGG+xBlRthq4H2LMt51jMIt4GJR+bfcvLCpQBs
h0t/Cxn50MkOrh+7mirLeX1KzHstIOLuQDlZ4ytXj4xZujyTn+PXgbJlsgjn4JLdj45yE7ySBs+L
0By+ysLE7zVYiKGUI+H8nWqsy4CjKtBP+lt8A56FsiRppZ+1MWuBPbmQY00lW+6h4hZLL7XbDrry
sAAMuDXZxIXqu48a9aNjfbkG8bLYtg6IzpWZRzVRK4ACuk+EFe4yR71tIWs6UM1yYJ2qkjWTk+WG
Vqr156JlLLB8RQXHgu3+4QeEyN0xHHsuyYyNkJ1UOS9dMdI/fL1ZvOOsCBHMsao08gAp9dawemdh
xr1Aaa2TdAYHzLydELlulahuoL4bb2gWPPesX6z2zLaamCEPnsWIR8Uk7XLRZJ+9cK0VuyLYDgOD
XE+6KrQj++QfFtwWEfzFoHpIikn5fGC6bd9zGOjoRLv32z1RO07kq5gSncH1m9P1e3p7S7qe+cp9
7aHM03ZKld+Djxq5Oxt2pGkq3/SQu9nY8y1RG0umaTE8sklVM1I44wvgUG8LkFywRU0kHbq4bhSY
TfADM0d38cqtoiuSNFMskk05ULXZWCSyv3Nbibr7biiWMJl4AUOKE3CGldFV4nIjKR5SOaueYu6v
+PkD2TA/7OYgqVs7dK9+5YRL5342PtD4FXrAqP/V6yQF1WdcNH5ZWSPKeKibtFy5wxf91kPlfqRJ
m0OgXhH6/s2iZXfAQcdasqoH6NtuGvYCkkAHUFkqKYf9OB6+sCmJ12AaiUCP4i2ZWK/VrvQWj0mt
4z5L0v0wMkl06PoJbVDzu7Z7O7LqJ2RWa9NwfR1baO3Fujt8Hcs44wuSVCKa8NCrvXpR75tnoJQK
T+dj66FqFjei6hCLfTXLI09HCWUHqBuijmVQUmSeXjK0hdiVpm2y9u/XZCmQnya14ucgsIKbdZ2E
BKAt0+ESl3U71tXA0O3KYIEt0AwyPCbI5vohK/HJv+q75u/3agjtMJzUPzGs311CPNjfQLK37HI3
hDTfPXWt4cbSl+CijT4pI0/jJtuPd8Pj7fxuOS6wrmC+U9/hKffGmi3wS6fojeEOOATycNhZKwN4
pKlVtTR7Tx0EQrjpQKGLldFSPxIC9LJ4hPdIrMtApaTz3dwvMhpF7cAGjWJCO65L0HRWkOef7quV
/W7m2xRzJ8RIJ4m7bBj7S/UIGGXUTwNQTmiK0IE3/mYgXZXUamwu11YTWbrUwsXdqv4rJ+Uojg08
1EQCjHdiBuSwfbMCx0eU4qyjpOaOxkhd4pV95oKm1xgTwXTvaXg7Pf+Y2RwN3MDDlq/XhbEcVw7Q
8bBuTEWa3sZ9wUfbUiHVKm/rj7P4zX44SbrA1EFbxt1jya77NRHbunNNq5wkDO95XktaQuy2rDKX
fYAFYTRudqFJ59ELo5vJfiQFhNepLN00dssVjtn3MFwRTmsHSh6WxHM3b+zkLp3Gqz/dMPmPOm/B
QW0eKdXfMI1+yg07CAeePAF7PS4QN0Jjz1FB7ftaz5mczdJlL0uu/NXXZSQu07QwkpNqK8UU+m/S
+ttm1szSOlMuweFmlYBENh9JF4S9OLcLC+Eqkt5inATLPPvuBLKl+Has5Vn2QWFEH8PijUEI4Aox
PcwrSNKFR11Nm/SUBQvLMJy5FhGfNtzx4HM4moJxoTuDz30rQ1gTHIXAO3rVfNmfEfWnVgX+Gyrg
UGtVeJ0+bYp3rNXf74n17sCwzTYBK4tvTcBbKpeg3RY38zu8dHAq7kh2BpS/dwHdFhnQzLILkcdb
CKZNgYHMHkzyOlddGlOMPdna1sbDdkqQ92MFUc6j5YWL/i36VYrVP4Dq3qU3j1ELzH+F7pMtSlAF
dxJ7C8fUUTVNSNL3QfvoDMmxsvZquKMFjN5yV0OcgRnj6kd2yvpfbHte44fQ6+AdvAmLZGInuBkB
Rdm/dBA0O868/rzNUjc4nZFhGYBcw51TIczSSwcLNg8TrQakWK3vjMZL/lysXJBBR8i36nT2s/bT
EU58fGANPJiINxk72ps+D/XNIKB+LAZw3F/oETAl9NNUbZPfc8Ran5ApieQrfvcQGtgRpOgY1TMh
V6nvBih82WzMXzNyim+JObMAYarOX5YFR944PQn42Sj2INypog32wK0mP5rh5gclodukS9Qbzh55
2yPOzWvoVShu4eZped51Djjc5IxXxT4WSIEpyoEeH2LGhvonCDwRbQ8FzGamXPD5M2EJA9z9CYNF
OLHYR71IMv+Mril84nuHEIIgZWKvRkNM/IsapyF6RjVGfoxTOeJXwkVAYDBPzpwqaewz/sZ+icVT
kpjZU68H9YcHqn/f4SMmO1l3GxCGj9/P+sPy1v7V60Tjg1jhdIOtUn7fD3ouJ1PlCTdVx366UXRs
VqBEqo452jrE1kyHxAqv76t3lxDnIOXZK9ICQ63q0Wv3ZhIDQJ8bZ0jfyToJYhK5pmNE7wzXLu3U
eGhTxPkHWkBdTTP6VPGiu0ZZR/rLaWtx1WfEp6Jh2J2M/dnIaCx0T8M8Gt3m/2uux0o/K2BdwDwi
ootQbsv1hHBsQ2KpBJE/0XB7rPQ+sLf1tZqKrm7xDWIsRGx4JDgaEEkpbuS2whWSuF2e4dYZByHJ
z2bvZes1Ibr0Jv8WYDGX5uTVlJYjqhG29tXpoLpUqOmBLmunLK8ZpavOMQ21PEfZVa0kyBN94Ssq
FguqQwDx+P2jmMTvEsbhEBJBummb5CjjKwCQozz0tFdOHGoD5GMjjilmMVFWJCNtlPn3De5prUA5
xpY+uFC5dUyIeN7GGXnqUM36cAvYJbKnRmIKYzZDeIfw0SO3QoOmZtWudbfJXg7XyTBDXg+wqZm5
mnstZvcxb+e5OLeo7HuQu1pUPulERPFpXdILdKNrCotMn1sK9C6qZMfeHwZzi8y+jaGZIG4dTC5R
ooKQODCyOdnDd3M26bij19lYWI87W8Zvq3NYhsRCq92Y7zmtZ/tIRCl2D3tUH9fj5UWhM9aOMEeY
z0Sv3A08qqlyR/vtvw4dpv+8oDvaTzRPb+0IvTHSZPlOl4SkDhyMKbyqOJZX/8DS7t6MzFyV+X8j
WI1EcdcIZ+V6zAh3dVoJQRKKjFgEwhVsZ5RkQEnzT071iWt4DthTYBg1CjRb5MMLk3cURp2w8PZn
dLG6v35idNnop0SyXicQL6utac3Kr7j3sjwY0540SRF4wNc2rtnKMCdgtxwigcd0FT8mVb8SXX+n
/4+s/4bP6prj5z47qjMeInGSZk8MbKktPEfJEYBsGP+Y4ongQUc7A0G6SxAvazNVTb97Ub1POlr/
QofOips7eifs1Fz/irvsp6iRsGysAcVa7w3T8M6cgfhOv1gnrrnE3qwa7286AmClm7B4gGEL/p0U
e04c6QW7/umqYJCHvMznGDaAZ/1IaYNaUkDKOj4MoDdqwscrvAV1tMEEC3q7vhpZLbq4Czd91Sms
psCdZKlWwod4sULMhKvPOHpORQHPn9gZ2mZ6i8Kp+l6XZvidC8zIYkDlWKn9C349jh9tE+N7PB4u
1mew9KvQO81qYIYLB36gOPlXzpDYx6LIoZRRxNr5PpvA31GcDIkfsxpA4dhq9L6KOxTisAPEAlzm
GKfJe8py0p3CvVFkiBpz3fpuroTxOyurRqHXNRznWwnE9/vlKAMj0mcWv48i+Ch0d22u++BH1J3X
j4WU2nYmBWG4Cwc6EwkK6jiHQA+4hqhTFF/rCcQ59cZ8htbl2zavx610l2TW3NWRHsKWDTeQKdPy
RZNPVTRAoa0mpMnjL5XG1Th9J25im6J3oynUxwES6bK/VFrpijNiT27eU9JRgVAjranRK4SOXKmT
zxFy9+7xVbj/WMLggLFuqiiLBMKhH3ATPNhS9qJ2176rwst3oVzO+o4KdSS4vL01wTUsJw4VgCjx
QqcEeqnqcmoeLYOe3SXv2L6xq1XcyteUzQV+eeRk6qo5hUSlnC/sLA8NZh/xhYOPKgjigzrqo0yq
ltpH1x4ryf2yMEFmM3Tx9dsSUiAdqIaoRHNjS6xJWNpNlX4fuK5SSgKZ8ShW86jbJU/gBgUor0p0
IYAcJkHiqbVtp/5OPYR7Qm87I4p6bpvy3nePAhum3IChV46f6jtBemkSAboVdX2IfdvgNk3B2CiQ
g+D7TOqsYXsDYrLw7+PHIrXwsCYbgdm92lo5Cj6JcoU4h2yoL5WAVbjwlErqO1zf3L6kIQ4h0Z9r
4oS2YiCPB0P6/XSeqbMvJQJsSlDLw8TuKLifQL+yTYLHbodUscEWRnU94ngpUnxntyTiCZA7tHGC
y7uFYa9Kpvinz/WhbQ84wQRUNdfrG64yC+k4bJ07Shzusb7UXfvLT8FWyd0CO06+NDSwEtbhTsEb
VsWMUxCh5cLL4ldCpLTIFiK6e9Dj0LDPJrUdG90BVaUGZb5NbjSbhFb8iIXx5XxalFE6XzS9rl2Z
YCjQFfG8/imbtJel4j0HSUjDnLgQOIlGSBqZuQG+otTUplWhq1sDqs9+lwa0ySXjDOz6YjGr0Kj9
OFyrZzNMmAmRCCjn0/eZaDAACp3tfjnRzysvampTRE9tCmQeY52wrFkyMW9tpG7pLzKRfFBBFEM5
dadGx5l4ZMc0gy1ZOkESdM8YDTQ4bfZ1c7GhTTZvzgeSdTEwLneO66DUP7Q7pTTRfgVgCeQxQgn7
OcbTLeJ0MR/7rfVZZvxAb1IBRT0zDnfyRfUmIx83P9NzPDcrmLJcCY1nu4x/NfxBdYrIRjGozyrm
y7xXfaKxLAw03wBlnGS/oU1V90Cc+WfCydPXPiKRByCcgW+03PQZDLxa64IMKp3dZ/fY8MfeqGGW
jILOgjNb9k6IO0zE0sbEcxyBwOG1Yh3a2TiZiiHUc3voWgX7a2GRXjokOWFFGh1OvTNqFkxm18wo
r7XaTaWtlUpw/icoPdlBjpjCpUMl3x07UaP9QqeFBr8rFii7bt0EZrYpM8EB46AE43lOSAK4UIgE
+Wwop+8IQ+MyeS0FSk/JMKOoyOqaS8WIQWSo0VZzDSArxXFXHTEmlf3C+OtpJHqgJEfus7QuVoRk
j1YFXVYwutgE8VPWz+yLjD8DUQFWj+zD1arZpwDEQuLm0MnAJWG8jfbZvanD7xwyU8V6iCTwkY2M
Rk0bzWyV/B3zA+1VUj44M5EYSIMbhP8pjegXUz841QTFqQVd1H1WPE/bxQ+A/hDAejX/VdomcBO3
2qSZjfBGhFBflWUe+l2e4PZAruLkP5HGCksknlaAu2jG/vrF7HaddP3seXccWt9dz91lmXE65RWD
pNUJPfKq8HtJUhE8glz9ddtM5k/fHiUFU9yoDL1zNtjMBYNUvcomMnilgMexx9MYHbsWNm/1QJ/h
QIHFELTFT/rGSdxCEzMb17Fd33RwKiHzQCYXOkob5QDufPrffqzjkxXwh3yEBUbof9NhR71KWnDe
FQbHJA0LWPZ2j/0I/TlYA2kvpgZ10URU+fEBGl3tZncDJ7SBPJy6ZmZ/ZqDPQvR3JE+RizwZuSSk
KhBpXWfvy4fmAizNyl/A2kvGdN+VxpiJnPJGQm5XaZQUUMa3u019q0wc0VOGxE54I5u6/Qd5/pPX
q3t2jrwjT6H3YzyeHkHNtR6XkFwOuk+iM1Wr8Wn3+hWgu4EcfKF/CjUppZbIwvoz1j/nk9ZJFAL2
g4lV3l+xIEKa9lucQ5BSEW88jObxjiNpkui3im+8gMqgwur7CW0sUm7PtZEf1UejRaY3O8Q0Uq4H
EKMuNlfiNa+kBcezwf1FjdGHpgn8clEFK7X3HVHXC8uM45kj1cnzeQrxBfMs6BtfnMVwj3ZDyqgN
Cd9feYQh5xRUbM+rKQ+jH6vCF9IuNuKBeL/yAAgStMPaclcU55cQMe7k37YkT0kKaLBUwtSPTVvS
Wg4CLEEMAd3hLBdq4V8I8GiWyFtLoR85KpWnuwwdupa+CSbgF5wlSAnQSkvvNS2EEKkFIfSU9m9m
Jr18wHZeZUtEGkKKbPY8CM1FqW3L8fdRSkhzfsGf61Lai+5DmaUySItJMmTzq0/rucCwbhbmE8xp
q//VtFrFX3nA9kAOYOFk/Q9DsQjx3p9BvxCUMXEbfH7+6NZBiA87NRvhCu8mkTH15C89HmA4QEcN
IhnGGsmYsUk+CvDJcBRSgCNkeKz5a0Oy3tJ33dG8e3GFNPcWEHFIE/ajEnlKM5UKfIhrR4T9Pwcq
oAX7urfQ+eBN91YDC34ogp9k/Reditjro++jvNSFSInu+bvI6+KCHWmdn//TSeaZNafIrOE6bfAP
Wiav1nYN7uV8/nO/jhmpdtOqXeDUekZPKn7133LtPybZ80OysJ7ISJ+6ECWrTJ4ST0eWgLDg8gHb
j11pFGYqYQWdNDIa1sh6+PgwWfHU++LFZ1qDidf7x1BgwRRQW8/+kLYXGQgpjnKd6dY2lKwdsYO7
IDHIHvwA0KDAw95UWZ3X4mV6tIRBro6QXECQ2s4aE21gSasBF3W6314GAvpImiTRuTTUXfZt2Xko
mIUSrAK9OcBt1Xipbf3ltTSRnIMWkQ+gXNENc1i+5x92dIvGSGwaXIiPcPJkn6XEmIrXBIbThm1J
uqy/UZi9LDP5Vb+d+agbhHVlZP2i4/vh/+gDiTr1QCoYfbLEAcPfcBMc2qoOIhwTf1bnH1Vufcem
pBb37gQ/Xw6E7kcoyz+eMW2sd51hm7tOLw98LLMjY5L6pquk8k/olEwjQCxGxQwTZftNpE6UUNQE
bHyJgwaHrQ37u9mbhXIs+Wz/qLdICSyLMzpTqXIe/G9hNH8Fyh2/YLzLyyqwOyrEMKZZPj1L9wyT
ZMrxu0TyAjeaorPdsGD0c2rxZ6ZTJZmDM0y8fkmuCkjaliZ7nNCuhub4pC6UtFiE9vCYzX11VJKw
NyPDegREAjVefef0XnQRfN9rWoyxd/dl8Ryt2wAjwREOQ2D94ES8ubCADO1wjQjtqkY/YC8K+75b
GOthiEYT/37+bjeszNn8ePTryPG9M8B0OZ5+0TlhhBchc/4QIjWnS0VCWLJ/YgSsSbAn3vJxGO6H
uhGiNDNeHdoAzJqI35Vkq7SqSuuaaX//36cDCBU+y/8jt5672aKHZKy/DO8juYMjLm6R8G9xrh6y
msOn6wl6wTPG/1CaAe77hkeBVOlCU8F4wjo+msLD7astd0uBVYrcINoy8lgKFrkspnA3ScOf2BcE
mRAdn8SArnO8VA7DRTrhmbrDRBH/PXE6eLrPEpOdkoZ3M45Tc7HmmbU0I18Z30oAA8cNupEdRv13
HOmoNmOxlN0ncdNvL1nKarJVkfCmmxEU2FFD66DFpc20KJbLSfcMQdm/etOnHR5OFqtWnaSR4XK3
2MpMU85v0ciXQ/tl6zh7gfrcFb8JZxwkXx+iaMBxHNdJQk9hivkTw8H9FDldaeRYvijhXiahYRdM
VI6Y6yOTyf4HxCFs8eiV2vM5XCUPiMEBA4HLg42NWJpMGmaLsI9gD8tzCbqoJRXKsrL0y87Z8Pfh
hXHVJcRTZ7NRBobRUP8Mi9wThqKPkXisBKWnrobXcI2PNg1PI+GfSaYb0q9uYfq6IBb+wGei4l21
FnAR+jtMJWSoEQGsVKWy3l9QMLJFjdeHCA8wcF9t2O5Iq6Q34erAMTAtA/AayLvtvHH+PbSQ4L+N
iMu4bNv7tZ9CPHGjr6VsU0P74BY6ZVcBp9lS9o3YgHdm9jClo/IdGuEDoLDK8gwswk+rzCFLGyqB
oOeIFWG93g78iE5++v2N1LiezCMRaa2I76v3W04hGfsIVjzEZa9YwIo4uFEEJKhAoYEkM0ghG11X
gpyNYKAlFH66fjG3b24ANxBMSZQIrnUqeHR/4mEWHx5/Dn6oQUNAssRrZlw4SUkPXZ7tQLXTqanh
Mc7tm3u26CIsPi9tpoK06sg5jzAcACZHX4dt3BtmHSeV2hfPLpxviNj3qGvG/xb831809N+C5/Wa
Hbi4bJvDwvqK7nv+gc++XB6y2AagNHTe97e6/AJeAfADVwhqWl8rEtucednW+JykdaVm4u0uK5t0
3xrE8Cf0gQAXAvz95BQT8HhomnTVfPh7uDzpSwAUSzkdqE6tnnMwgzf3333uKVE2r2cEgzvDkczI
kOWAb+R2rw/Fi+Jt1fpsOTHbSZ77enFvsV6f1Dvinh5Iqv0o/jL/HVaV+FExKe0ypl7EW83rMv+U
JPjJncaLPsdpyeVESPa+zuxBSiSD755236qx9bjpHDaHsIGEzs+T9eDm7pXhwxFnsAUfL26Vh+0h
Rt7QsYQtgJJUNGM2azfmEQdIQ9sC1LkXtRz53tX+sjuF36iIZMY+x2zgqWgEfkfV4eUk9RK+xz8z
ze/md056eDZ1M1BAIxOGVbNfPZwmN6o0XlUNq6wZCuFn//LsltKwMP/tRrbfdz46CYRdwnJcXnGD
c1kMdOSdlhabQbyKFjpoVFedRHESkupu1EEhwaN6kXdibDXHx39bXSAA9owFzN/fEwcsCrlvvY2R
Y5/EUfEdG1lGlt5BkazFon5/89rlpRCqUiGgQxJOzyGrr7s4yEY62vPPgQIxU7m8NgEL0JdZhaUN
SW0TgH4wvs3H63zv3N8szOOfsMb5KOFZIVxAZZWAsqSccuOYKl1MstVAAOA/R1aQYX1+MDSuAzqW
TEldR3G7Uq9wUbT/4o/0t+fVs+N+06u7Ep5Dcx3x9bFGIO0yfm+MbcF2GS4Expba+Tv8dsYieEbs
xjU2Bo3xaGSP/sVRqaeC3t0hf7xLqUkbeF29C2fkaf1dKveatRIKxdXxzp2q30hRwadCv2TFgmfM
OnaqDfIb3BQwiO8F6x5Tw5pBkwx/7rL2Vy4kE/VjMS25JJXhwKHSfvqbW6UWdkg2pJlD9zE/ED5r
mkm36jbui2m5RMqO1pTtA1nh9jraEW2s8sGRkE9akwCtqhsX9vQ9r7lH74IobHpqd8eEvHSBxecs
ixURadS4CfnLYejipRUEXt7d2mW/WKjSq8lhOQ84c81GAZDnu0nF7jCN0KACXveoiG+oi8/ncWtD
hRAkBs7Dm1FUGxU3APiyWl/P/hmtQjpLkUmk03C9jJb+FT3orFaF1Rx5cAedfPaxa1dBigL/+/f0
N/lirdMzFY7hvBN1RnXYwIqPVUPtamoZnzTCQFwlHeGQ4UgqD01r7RVi0cf9IdpWCCWqz+y0Xq6U
cg1rn3P81OJvOv15EIk5zaqjmUf2cE80Ao0B2qfNxCD5LJt0tLDam6Nwufx01WetXNAFwsvizAQa
Yv0H1iFhAlG9yM61830uXSjAnYM1ch7YYZm5nWAE610yoCV2uKUCbZTXFtKpYMXpLdURxWONfyh5
uIS3gz4PW45dg/4kJHcx+C7N3pTRQN/v4dpazur1McDEPC4tf9RefAWey7deRlhUKRjoNqEjqqns
eJlZvqP1lGmWDygy0g8jw2KF0XdN2/58V3TM8MVgBKi7ImqIjPfPKxuHhA4qOHRL+KQc2ffxlSpT
V3kGCHUnx3jHeJMgOG9CIfkTI7KhfT0dTIOMu0jI/QVtiT0UDIoZ1cxih+YhrJ9xI9Ae0kg5xyrm
ALXmhJ7go8OFxVs+D124+08DJbTGVuJid4I2IQEsHpgDxT3s8jGR9am9dBV8JXtEANMsukN9VGUo
R4B1CCZxz0qSdK69eTsNMn6WlSUaFT814P++QOarW+4b3x3iAINZktUCpVifdF/B7loxwOEqcq81
jf1Cg/4Z+tLEKd5WXLG/Gn+xKwXy1z53lYAeeeILL7K8qw3UF3lv9ODREo0nO/6h2d2mWTa9A7ZE
Y9UlvELDmjZfK+WqjclQHXBkN0pTGQKF7oEP/m3CKTmzG6EGk479FkC2gOKFkCOYfMhRDAg2LkoS
+YiUhIM4+1DJXd7b+oi/IRjz/cs5VAp1QAzuWQfPULCdlqT56wrQQzz5I2W7hNVOhCDhQHTa2xHx
7m9UyEUlnBPXAnOh3c1pvG9crE1yPTdFI4Afr0LrCa9b76LgtiuY+r3/F/AC40rzCOIUVVLkuRra
cRjMdbvolICD3RDZt0oNgJXQ7cvaPwqD6zxbKxSg5cyIFWqTuFSgwvlYz5Qu+6DjNxJ4sDSaKMbk
jpJafxly6q30gQa0AbPMS7czepY1u4tTNpO4LfRjPdSS2sdfP/ZjZXR5AoyNHS22BEXBnS5lfSHJ
9wWPMjB60eEbrFdt64PIp93i2V2YGvHJVyc4QYUyBQHTVnLLu3+FUU1jICi8f6OZcgUjy9AYLiPo
w6D8wfNgQhYN/dd4wP63My2HHio4cgg8T77LPNqKESHfUn4C0kWqGDYIun7ig/2Ft1wOY/WelvxB
LwU5N8tdsVGhIX7t9iwnbKAyQ3YIMbBfzY/ouES7AQPy7wV3AQ6MY6UdlnvHILTR3IT4r8LXcDMc
9t9aoKhAZaOVKvy3Abz9ay7oZtnXm605d4pnFyCUTHZOKAck3ZTYTgxes52+Y5LqCShT0/MasqbA
TzZDf1Zfmg4EpF2uEsKRc8leyKILt+oK+5XqVp9h0Kd4QIP4+mCnmXt1rjDxudK+bzOxY+g3mjzi
mUONvt4V52uJe8xHkRpG8oh+xJitIqzeAHusM9wduh9apqrZTZ081vXAsa+hYLQJUlXVy6Jo6fv+
JDwNerNS+j2HVVeOH7aceFu5LL5xgufHz1Q+c8nIzYmQ9PD0Q7Qd7faCMrpk6SPEzIuwd0ATaVDP
zc+T+op0NWeq6Idpny/mv9RlBHzX1zZlwY/IMu67AFQET9a+FJy86JSCFM1N1bilQ5RES4MIV386
Ecv6hJJA6Dl0oFGPv8lzMPbzOJl6J6GpP0R8aJL15WOHkvmchK5nScS87TpbmZkgQXhleLEy2KV7
ZGzho5Q+dtY1toB4XtV1XPm37zVkA2G+HhucgmIWqjkfj+zhjC3UhrEvjmeT3wrHWXropDx4c3ZP
PCLkyrFeHEJ4dAw0VA2E97t5GMhxt5nKqGcD4LYC75AX4f7SNGU5ktXXGru+yrr7tHkuidy1IEqN
H4QqI6ugsViWpF2XRr0kZYuro2tkYiahwP0Uz1p9O45d0goqDsH+xGuYxBiGfZk7KrKKB9KXpS8n
wVl3YdsD4JQEQCCobGewDCRfSa1HmZN5CtEmaKuOw8mcJx5wRUuETsQ60NAfTCxKGlZ2Qx0nP2hZ
5ObgZO9BUcpt7BozPl0ta4HiescI1er/66QP0/WN14qZKMI6MdbZP9gxOajwPF1EeOTf9Zu9WcRc
ugRkBt368OfkLEcfflM85IhEwe9opT9Cj/pd5Hm+pRi6/XlXLROGWRD3ifjq3Gc1wkGFdTBb1opj
7MEJsbHVU53+7gTdZSSq4f3RAMy6+4L/T2mD2al1bDnX/ESYXn9OD4IGf3Y9MZfRubTcFj0+H1Xh
gMoKvkCWMVV64sFw23uQdz/aFM8P4DatdkjOJg/ljhU6PnYL6n97bgvKVL22h1FU6m83YEq+c+6p
fktw7foiaBTEoQuzLJArZJy2FUIVHSHNa/TPjKXOMMK0GNHs6uFkgnN+dsJETZbdyUz/tOOaDFSo
BUuWKIkTiA4obeB4m+UDJFNX49D0ZSo2ewWNTs2zW1/DrHbfIIGkXNkJProEqkoniWgKUQ5h+8UE
FNrIADNum99jWRFKVFZqHRVUcfwwb0vNf2ZZj+Z0t6HL+rpcQEPJOE9QnOy1FufUwWvnfENf2ky6
W/l4M7DlbGqsxzHXQMmnCnDVCjP35gBGAxE200jAEO2l6ny22cq+S965etPgk+/D4gXyH16T5f2r
SFAAevysiyddc6U4DsffgAJidP1tMR2NYgDXgdd3yNiz3y7wkt7B/oBtPgqn5FHhMLvyBZQQnnau
Y+93ObwhGvBBNDm57Ybmf7moFEaQdAODWQ7d/rklHie05zbNJOW61yOZUd1fJDdFyEhwMKUrDX7C
lV1wZYVPWDWHMGEoNg4GrNqcBZTmMRsrQy174Qmy9qgAqPkHJPL28CqDHobbmXsz/x5D8XAVHK3d
kDk6yDmDxMprBfYQCgWykEaAm6dogfSI1ewsYeGkDPUDF8S9GkyOGh1uZMnKlufjklyIwglWgtVQ
3qHShrG1twS9w3KUQgivx5WHy5sAE5kbPFHIOKMKBQGAj1cQ5d2rd1TVgq3pq4DsZT396O3zrth9
Th1maivySUz5i8jZ+TQIDje+EfJhHiSAw4r2p0OmLhlPURq4vwEVWWuGuBQtvOaErM8JdxuHwD+j
2lnV6FvXkWBn9oYF3YiHrPjr8RsqJ6y3QduPS/kju+ePoKK6LXFV4wFEIZ38UibTtcXC0hynXFDF
Y8NJDNjNj/FWlmZFQjU6CqNNaFDm+HS9R/PoxgRjspR3VT+/79RYp4W13PqrdAzETJ++QlrWQbgo
wKeRiaA5g5oyS0vPrZ4S0hLrlDu5JU//YZdyWmJkdow/6OOsaOzX67W0x0bKGOevzcB0rofyT1hN
e5EvphisNbLEOxhMjLKq2b7gYbslPfRlWzs8lA2oZnthPDFeT+Sv5KeXof1bJl5VsMFXDRs5hayq
93h/ZgT0p1q2CP+dw5Q8jxYiWDXaKxgNi9knGi+QKEbaP3xmntJYBg4VMh6cfNfkM+urndb5JDTY
8bA4I5XA866P1+FKLFEgoRlKgm6NSp9Lb9XYl7+i8qk1jzqcoKWxf317w2VmxIX9KBIKSCZHDmiZ
dzATKqvzmnv2tLtgkafeITiTnhboqk1HM4sHAH7f9PfRrPaOGvfHed8qbgFHC31l59QPCV8Kwi0H
8r4imhGr7NyjacrODCQsD1L9v1bElNnkqFPxO92W3qXQoQG3I/d1fV8eVyNmWFVN2ihoofWMHVYz
1ioW/kUTuWrpLs5LbSAe8soOyGneNDE1wJUTrPPpixhGRZmoyxc9QgaVMg27KAnlwZ6WsuDalBKa
PIeD1ZPs9ZvZ/DEpVSLHE1UzbCzf+0kD4OisK/cFbhhQMqygxHvqHs1Dn11jCV53W2+sn33r0XmW
QSJggTo2mpoIWqJAR5IQalZMrbYq/q4tM4kJutPXDOTmMPH89lm91o7vTrRHMjEzjeB7obKPF8mX
H0putvPIhg7DMgpcPtODbdsruuukPEyAo6k1liPL1WzjfB68FyrZNryBVmraCjsU+5WebmQp0l5N
66CjL+NngwU3AkuYLbBkJGpwy7E13GD7rkTjeYMIbnOKq3W2f1T/c7+fy+Cl1SNltWDhwBGplSfb
fv02wuvhyoMmOBnt6bquwBnL7i4m/EqxByaAph43Yu+a3oug2Z1w8je5pKeSuDb+bb0xrjBOOB9n
YbZhFOncA0TQk2DFQDjEQ2dwhBaNDpKwdHq1mMHGFsYFmyTc4OI0cXQRmhr4xDmG/3h+Kjgzk1Vs
M8CVK5PDBYRcgCLy/CMOAd9YOBDrTGvQguDsanBOCXXzQYhd1Imh5D1H0Ml+uQWPy7LggoUa5LBg
Y+qRgnt9oJPnM2CTW9VO7MKw+T1afBYHarRfhnqjUWaWASudk7cGuu2C5VC0WuLaqt7uoI5Llc2N
P6iWgxJ4Zyhp1TeNfbQFQjtEXcETq6OSp4tG1DRZceG8OwqOIKEbra96bvSo4e9iV7qQ1YmN+tnP
XQxiq+SzQX5vZ5nGzzxXrzyPSzO3hc2lal2zqqnMowdD7vAPCgQREENujVb1eS/n7ETy5UJKSJJu
qpT8DvMFlELi5UQO6Kg4Vdet3kmdnVh2FzyGbG3Gcc6qytnYP9m2qs+DWXHz07a2gUvxoFXVZAGV
P+6iVikLjmc1DpH9kaqYQC7UxRnN2N1Z+VFQn1SmqP2z0UtRPu/IkJHKgq+Ec8y3uptMaMIWdIrp
uOV4cmq4M8gZzX6/5e/PzKhCIHp0O0JEJwUTiJjYTYFA1rQZPUrjVJkZ3boj/eDFremkhsdX+Qyq
kiGMphmnatNALdS3pyJChReJVpcAQOnfZ4pQvrJpd68D+fxvwNYU1Br6QlxoGm6lHrHz0DB6Nj4X
fUHapu86M4GkFz19RGwMpNa64+JYfHA4dKliBKk86SxWWOWmbEtm9dtp3yeX7luUW+Gkp5176egR
tx4DBZ0nBSPZRDxq3yu+kIg29n/+000HErtuzkSpH7fZzNgln0TmjS8NLhhAxUFBGI/GCn4YNsTN
1q7S4ForUlWnO1rfOru8RPlbBVs3Jqb0tYwYY/ISBMSpjIHiUvCRiYstQDz8l0RHyhA2csv65wyw
hjjGgFT4Aglk1v/5jgZRvn+iM+sG7DaW/dAux4wsB5p3IPvxycBczbKMWhW0OUPqjQRm1Gw44Uei
gfT12qWiq1CqYy8sZ/w1WfWRcRDhRmlw9mmcD+lPViaU5H9/z8kwaVTPvGY1vOZ4Zavak5dbLJMv
hj2yHDx+AaDoHMmk7KsNh6642JwUrT1ce6Urzu2VExqSwQRGHo65FavB3h4iesQb82ixWPbQTxBH
/371xb1lLK3i1v/e7lMbkcWYKyLK7iR6PGPi5oHA7FmKVJ7LIuWYq5V9vAqdWJEYkLcKBq+7kUrS
ssGntwiG2PBp7UTboPGoVpCMnujXoQ20JsFmljDN7rjDY38j/iOnhrjY2lgAQLZ/Ht9/xWcvbyh5
nXaU4HQqCl/KzEPx11+EafxJeTfNG5bRuZE+TeE0f3ZXfRWkqFNP9wdAE2TVXnOfmL49EajR2PJ0
/NCZiDes1k7m5Snejuq/ArrLvHn0mpBcaPNMUfChVvbfmqWlsMM1afjDg6jTXpASGeZOb1Dcokpc
fpgZNSUxcOemKnJzzHtNOPpv7HqF8IurLsj5TIeWRXImcYKiRr5ukkt6dJiU1BrEIVJjqjLcE77k
EQ7Kjg/XiIGRdLmzc0NyU5UwX3QHlWMRFiO+qvrVflM735BQ5fk5CwDsgYQlByVvAmxS7j3/6wSX
YpsZt7o8uo397fFcxDCDmaGHE66owjibB9ukz7P/1p1pKL0gLPjI10lukuB5VcscooYfW7wzrjXk
apUgkdLSqP9yp4IpDx4hikzRrQNtcsXhmTN9/bNrlqUo8tnLUZ7reIpItSzED0gZTKubaizpYKFy
ZKAMukqckPab8i2UUDLS200np4wAyZ+wl7Uh6OToXC8+BsW2Aebm3cJCw1DLmMpfkS3tIp1BJo7D
mTwlX8LL/H9n192H7D8hkrcfe3L//n4rWgbbtUsr2IOqUTCcl5TSXShAqfg0oPGCPS3p24WkdsQp
OT7Orl+WPRMsZPnYoZbMjMp23WJjPUd+++GgbL8hfDcNIU3Tn5IRIxWdqZdD3BcpwFqGC+veBWiW
sVg0DNTb/Eq60Rc+OjBx5612E3dB4YAxbO4XNTFj0vO7sO/HrIrT+G+jnk5SZStoKVtVi/TKcDYU
AR9jr5PSCvve5zma2FxMIXSuTE6oDUiAv1czVlGP0EigEd72XhBLhTzKS6JHyKb/PEsDAmZvSvNN
F3IYtQqtCnA7ioswZqoSU6bQayqXNLIuz/12fyfKLhvJeXlTllVnZFiPgjNvxqxV8wITvwF3MYe1
F9ju2RjD/JU6s1Up/F9A2EhX2wg2LU8Jk51j6+n1zwCAmCnTZr5RlIMioBV2+/GwRJhh8gygCBFk
IJntp46hiOZ4C30Y4kRcyMDdyKNj2JCdkhq/MO63tVukX2SbwgXcDMTuZ3MJRMu5hO6fWqkY30tb
R42FaJ8zwmmH39cwqqt+LJZJoRCtCp3xoWvpcSowAfgxmw6fiAZvvExM7tLKzJX8cG2H7tkgve13
etyoxMh3oVDKnrsZpKiEc47FSl1/OmDVsT4/YG4LeN8ES+MINmV4cTC/kfsUkm8E0uPCINYPVhxU
p8EwQ9ZEGlXWi+7CQ2pu/vWpmES7ZXJJyAfO8KE0f/06IzrJs2TAYFpaWssi4rQRu43DTm9qkC7l
1m3MFGxYy97sWFvHmZH94K3RVs3y1Hlfs/f/zPXI/Kbx2jWYdwvpK6Ej5i1jx3WhG+vjGHQF1ZDY
mMf6CWQ8+t9DQKOMqcn8h5LY8uiYhNnrALXjkWm9jdYlvpXaBxym5GQEfW8Xmoe7pSl9BV29s4Zz
9hN5PY8hmE46pqVklDX5mgltp89IxQmj+KGYqkdsVVx/C/i4HlriFpLjShgnYPS7uA6+tqukiqyq
0vymDZaojWE/Va7vBHZ9g3m9V56wXdErZ1bBU4X6NBMxKbCfoYQSgReWz66nKq2FKq1RsNEYdNk3
h9C9JtLSVrYpt1Pgq2kicLChXkoSc6kVwS5nN0ivxgaZS55/OKvIK1v+4FXM44g+6JvJibvXQRGR
UnQQNPl/Uejk0UrWSfHXLX2iMLPOz7rnmJU0HsGOjjynHio1BrO8oltYjyEXumD0k8fmRnEmZm3g
uTuvEyoFc2B885xG1/y/Pcn+hfHLU3pbdNGR2g3UZ9/Idkha/VILOp5XF9rfnEYcTJmAsJmeZScZ
JIzovHfdEodVJf183tyg9mJW+SNtGJ/uyjakXOjdNku4HYt06zLOhX56w9an7LnUhlBAZ6PMyYWj
xaOCsEBQjQH+tlRMX+ZjRlUakKkpSqGT1TWo02Zs7BLN7ZKUr76L6rxrpahEQV+9bS9imiU5ZqVd
K4mmOqZKq/Yuf70T7WfIjx4Ke1wPoaoF/bsa9kDESjbjro9S+cMpjyWUrdXsL2h3Qs9yiuduqYEq
nfEIYrp+NcWyxi9hUXaeB4Qw1P/U9uHdpzHjUqffI/2Z1g0TfXTvALVAqWzFV3B+x/P33t6KBYG0
xh72m7ad0Di9r2j6xCZmhs2dbwmWGNUm9JMYZhDeEtllFu7waFL6o0jbmobmI5ofijKd3IdUlxax
+SjhFsbaSpGuNAS3HZNQxIFDaOKk2hG2627Yh7MoJ8MtzaERLwyfF3whjGoII9ddB2rlTMMbbFna
VpZ5leMi6PQG6pyvZHdlJDf9JOETfnJXLatdFtkizXVAlhWBtOHuMg+T8L/3wPtp1hs0lRkUaUr/
HuVc1pkhF/zrb2v15V5jlsS5aTReZYQsZ4AoR4h5AR5R9/qMz86zALr0cB45XyoTNXXxHYIRgMas
TDwUa2ND1Nhp6Sfda67gw2EsX1LLHUiYX78XENaeeTZF2tSAH0f6wdEOE5brCyQMbUqPBjadqLgK
dMDYygrDVVt5/F6h1A7K8Cdvr0gb4ukucac44FoXOh2cOAgwTVCIbdOGyhwZ1Y6cjPbxqutkksLY
KJahlI7IXSZ2ciN9nHPpLYSArUGCuwzNRFsNBrdLp76VqyXvRfp+OtrkZMEgfNYx3liKuOucNkol
15+71t+Grnv8PsN8+J12K1IiketW3Iy29ISmMOJf8ShQJzfCwOOhgE3HLj/o/hj7zqwb7pylk4wZ
qfZjAxQaQ5SZNH+bVAtN1jESRNsYf3HnahVF6yuk5w4wT2kdjZezaeFIgPoEf3bRZGVYms4S4Nny
59cQ0r1Ue4/AdTrB0GZS1hZKU5CcWmvQsfOCNDM7lD9gUXcqu0V0tWzhcU0AHsWeSsvZdpbvkcvg
YkQn52ZCW0gA0XfUarYU+BSeQjnJrWhLi9Cgxi+ySBb6iIzpCH6QIZFxXjDzSTgFe//P5DBxuiF2
UtqeCd6FTfIGNQdcoTzwIaHQ9bqd1j4TeidaWy4L8MTv2Umq240eSTNujUV4nk9eUef7Z/Oc16VN
N+KaE1RtALpJxKS/5yM9dzUSe5mvH7EZJFlHM4xm/lmK2L6VC7rp+zKqCQpnK3lnHre8S+qVCwf9
4uejLUm7hGsTOBacTy8kzDk3tZbiXxWcfEbrdiENH0+4QSBjbY3SirmNZgo59XuIZEDL8pvTlJg6
qwckpaRSucF37gGxcLJW0ji9J+OJyxsFHkQ7mayPtIcbwfA7R9NthRjxv5OKuOXnM2ZD0Pot5FVy
Qs1LRNYDTRTpEOnHIMjKtqJ4fQjOZLuZgkVZEtM6lc4CamjIvw+wq63DXagyvW/V5cD+w/uRUIy6
U7hPYhQ/Zg/8Ez1Zp27duZeahmFeYz6jmXBgdr3fGu6uaH2bphXYtPaa2NVlK2OggHdwhjp9hrg+
MmuXTgNFn9c8iadb4w33cRcjE94kdAtG8DHMUkMveZvC/IotEN82RU9LCUJKPsExnbO8FAw828ml
WYcWdZ62GRHVrHGqcay/EuXyyaz+UbrIJbeEn3q4zfeiFrPDii8bccNoC3NQ3OS7iA/OEANytGuS
+cCLocWwJOhGDN1vHRSyf55GhfKPDdVoGDnWak2P3z8oz/gb5wdXxB+AglDSntOPvqkKDzMnzon2
qFMzd1jLUMgHJC0Z9T889nxXPfHHZuH02kOvVa9n1HR43Ig2TWbPsB2ebPgL4fwF2VDE97MFXXkL
8nQG1drk7y3KpgBqUPb59GAoahbkzYDSgWHiZDXxfMQdcEuQ1pOOQo6MHldnL1jUNdnjFEfQinJb
3yyajojV9RfhzB0X8cEEEZ7LCJK23RsOzMMAatsWnx8Uos39oHS8TSBu+31VPs4rb8l3lB+Ma5f2
668tuUdh1adAgb/obfrCFrCtpw+9TKS8uHmMho7cZEhVTtBy9RVGVmdL9qs31Lx5iEUGDlcN50+r
hjDlod1YLY4H0GYn8jeljPRr3qzwiU+Zi2JDmCDeZLErvXAGmSxGrFMJCN23tmEoScvqAIzEf0Xu
Se2pTlZ1zZ9CR/+G6onT6SRAXFFmF7Yr9K380dZ6+tvtSivFUwElpjhsa0rRHi1qIiY0Rhf1O9Gp
WHYm1q+rJJE6NoTiZGi4uGh7bqs1x7+b9hT0hn2DAw4vBJYd4AGKsmyHet/6G1OX2ZPi+Xw1E2FW
eEqYt1OHh5OnV2YlW8Q9apTDkH4vFU72lJcd+Zkprus+1BarLSRxkARyNGxIfhRc5NB6KiKyzmZo
pq8zjqvj/eQxU3r/2yEi/2I4GRDaoZaavdcrR/BheGOt11uOCkCezBSpF/1fz1ljDlGLiPTdAl1W
I9+A4TOj20knFXCXLFwRQkJX7oNPeIqvtlgW18Xvh/qT4Rg8UhV7mjejCVPA4WSHbTuludyb9JbX
/tKFMWePO+0c+8r9mL3uuAW+KoDfQomjLuKwikPXt2P2LKcB3FlvlJzgVBQ/PzsbjKDBzlPSUYVn
qTrYIhP7UxhBEGn8wUWon6Dozah3VLYDo07HM9RN5sj3/z5qLcnFTdWiG9CJPFLDQrsCrxHmDoZo
jF4w2KWe28U8p09zfE+/MceGQ9RfTf069PR4sU5zzrOjHPa7Fs48AS2QW9hLLGulYjPaGl6nhEZ+
qqVx7CePIgV4YFQkAoYYo7YMXN+RIBGpfSFS+OBRFsJv9UOht1yIjr9oNviak8hqJ3hl638Ii4ga
DmH1cI4+v1khGg9XqBa0Ei9Zd80uycM6Xm625/K0DV0Fj7MjKyNNhJo3btVqsK0RPUkMhRUA7BQQ
lS7qHVe4u7kAbKcUysb+b3/cSVq2AYTtde4kgITFCmPxEk00gbzSN9xII1QO2lv6LTSy0Z3bcw5I
4dMlSWQq+k8IZo7foXCTxWqCyTM2eGGo67PP+XKBVo/pCOY4Dd8Y6Tuk8zgL0BvpKoYViHasa0h9
OAAfoVFWg87MVTwuxp/bEd0yYvnMaoSEDN2b0yamNrQSnPRHHY/WuLFikNQqjLlg5P5JLGwCQiu1
vTmmmKW78/BF+/b6eFxuLBvDufUusEGtKhj/aEAMQAwYY/FrlDuMFuPkTwdxIxBsUvw1OWMKElA8
csO5g8JGlEa4aWeAfeEXJjUdpuNnaJxBn3UgU8BiFzCsl4rUpEsv/I7uTQgLLFg2KCAXjZOLG3Z1
5aIZsYi6p0UCgHM6baeulBAAIOi3hnA4pjt4zaLmaVwY0LRpqfZz8d7/pKSF9jbyEiA4eaa4MJAY
suEBNXuWrpYse6QDyPPgIDwqVrRV2fROxb2JANyXUdQCta34F4Q01hYS6/ODfjTpZN3zdMcU4ifo
VPgfnCzsigPbPhGkM3pxJ7dCV75HN0+6dTnX9eH4a4h30pJiBjTbzISTo50EufyeG78y8nmlDY29
iOXSZEDHDVbmTLYD7yPj3JmZZBq9cd9R+YEMjA8/ulgc42jN3lol5+tBHJ/Nbzboogl0VRUFkshT
pNxRscsnU8C7LZzT57MuxRsd5+w3Bfn1c3K3n+XZVw+oY6Nh9Zt5ENpZnlWCCdefBmfmUFfG30XF
8ZhHlnlShFOzN7QYBUx9jU5yqU0hSxczPSJh2Tgve44dIm+lzmHfp927E7yV+TkEh+2IR4wY+vkI
JMFiGjlvyAUYVJsmH94RNzMVXWi+aCkm4p4dPlMn8s6v6ZzkdnxsiqoBccxYesiulJRac5fQC+qL
dkuDpPY3qT0ob9/w4jZoSvSo77Chin2Oumy+5fgxfvgj3NEYsFnz+IbDmfWpKLAHk0TQSyL/hfjg
Gk2qRwCgOwVPxi84e4v3VwL7jFw08IQDTse/CWrGyaxaQZq5gQRRa3YHionhpYv+xlPB1ERTuyaF
L6X6X9+qMYOVqAvg+QAWvDDKzV6xtM+uAE/pss5wZg5fPU3DyORqSUk4SUKlT5k6veQidR34KebR
Xme9ZcFzYjMcaqpcnWKmG/FRHp4j08ZfWmJn/U8QHpD106Q064St9SoC//PYdeevDyEGTTf2p1fY
mJPiGDNvpwtNwoXdnX9tNKcBeH4CgKyek/uZJVHSWpdFc2jU6AOZddbTuIzJCEKyhIqSEm2BrMPz
vpBJbNFfFI2Idzkxf95sy3m949/fC6vHyYhpxDCyXJagkkmlKBIlVNPug9oonrbBvBRY7HFFgsms
JIpB/JHGyp8+qnDxEdMd1Sk9z1ea2fp/2pzuWej4BI2uaJ9EN2uG3xCb/cmpjrHSHaYBwR0ltmaS
QQvkhWn/DtX+gBbsJnAIUAQLGLaSlJQm6eba6gLbSUHipfdOnSeVwpJyol26zcdheMBMb7r6AqTP
nuOpCx0nIk1wMOjPOVk+koYvEKSe43VHkzW4313a/CR0U0l9QUASkCWUg8sRpcRkjMVCbHIHFsuv
dYH70EvGp+p7YXQhsOncvj1QSQsw8bmhmtcUhjsc/UGHTjn+8Ipvnq6tUsJNGm3lVlkJf4gSouyS
Yq2Y5Lfu1v0Jgo+Qz9CFZctmYzJHPsPCmwmCG4R9tNevwi1DWOuL97BwMLbieL0XrphQmBD5IVu0
b+M8Yf577WwveIxPfsF0QpnwWCJN7bQLNNyo5Y7v/RJahho+eXPfSHJh5A2CdWhYoQ/RXBluu1pB
mxjjOQf3z+TkvxDdXE2zNbQ/JP2/+WBZrtNHSj7Ms9KUimYWViK1lMNx8O7INbHafAylp+t4GnDp
Cnqmmr+BjtwU+7QDU5bKmny4BTeu9oSddpTBvSPZ5xorXV78PGrUMihROP5gxEspq9HMbbpkfwHo
xQTqPdw9FAO9UzjLmcMSwMnLshqMm9nX+q0WR9cvJeJNqswJRA2OfE8BHcNx9ZHquszcyD0LqPtF
8KGQ0gIQaNi0nIWTzc16XQTOt7EvkoeUA+63SAM465uL4IYp+DHDn431pYBRGCjptoY6ClTE1gJ4
var2HTy5yjQHZKiDNa5SGvTXvhSAFCskkveTPTzxyTXsITdmnKNYO7gev6YKL6TDzwMsYnd2G8fz
ra1VTQOzb962cPcgQvVyqP0QdCqNWweKSzbwO/tr+ufW/OjRuzGqbW+/bYtdDK8GzafVKKLOFTd7
60IxHXUUyBFIgWvrF8cVA2kN1rsuPdliLf1QVAGOiyiwsXkt4jWvFhx3g8IlSKF28mUvBsslhoDF
7pQZD9x6XNzr1UvBhz2VZ58FcxuUjGqfX5jEYuGLfLwyJgB0ji+E0MhicxOOE3SezL59jbw2c57z
ZS0O0u3SjLbc5kIZ/B2kDVZ34gGGuJoPja/10JuwGgDZhoYqlr2Cu4gr5r1MRHn3XxFLH9cgi/JG
99pPSIw3fn1C7CFR1UDzLvhJXTjVHM9FY6T1RzbSli3/iYn9Z04U4elvQJnbrZI9mFFNG0FspCvu
LGEFXaWe05PDy81JlsDZW+wiNf2INamtjnAorjhe1hYn+1/+zIxQHmoUAhOQW8YWiaYnPiZQ7bBN
Y/VoA2zIuP/Y2990sSE9T04zAhq5Wm/AC3N4qzmLQIzkwaxiWwkkSGwMtiBk9w6g0/8cSZu5Rj8x
NHFCWh07m9gjcyzfJAc1ZfAN2b7Qmrtt1dhHm+6R0XkJ7JH0Y5gweBplaIDzmyyidQ+bTgj1+Ogz
oLpf/XUPbEfzcOF96QaSgSdx9UFTG7YPWGaQ8oBFSpXBHT8qiMZvoB0PNximBDTpVvFHaygs8+d3
j3erRwPiZnQP9Olr3+armAibexp/Qq0PiIk0nfAXhs8ErphEB+Gxukaz80zXGKfJv3vuWdLECF5V
faqdUB/r4EafybAolOKDW9Hf35JS5ocuSWgsDC9BYxgwCaeeRa9Uf+xGAZUiHgXvdYJwX/K8af9h
RrxyCkewmImGB2xPZV1UTrHa1RjVGBbWNotFP1KASv2ac0deDDLo7J7OrC8FeVXb5AumprWGK9rp
CjE2BEZakY7t4G1PBJLRb/Z3uk4S2X5uisaqvoDsnDFPhqPFlGoJ2uiJTXsWdHNsCRjoPZuFr9o+
0ETaW+ipupMwXxYHHsTEpKBo1q9mmOJ1dUP+R231W/6twCsbbYXeZm+aY/YI/giaHS6zRpW09Un9
h1zfnEKIKSXFPdmIWguoZvXFir+2w9rM9xIcboGhu+qoCwVpvFCPdx2OiBVjQPvjsMpE6pLXDgEO
jdqOXdbL6nkYEefJVKmNUcoLDwJ/4P3G7L621xYyq28nlsISNkxXrfnvvTm2y4aFE2aSxr7m1mkF
dAwf0ts26+dPGyoS2TCbAgV5kLrFQPDxLpooPLgQQI/Jk8c8e28FPW/C6vbtWcTLrqIok6yWH34w
l4QA7lYFBxk0c8d1mMXUU3fB1iI4HnrgBDRS81ua2OTM+sZLVBhTt/5Es2VgUTV81zmPEo08LXKn
Pd0UIeMEPFx3qBk6e/ygFy2SqO3nW+w5qqhoiiguNvAShx9pbb2DtQjm1Qu3UfGkYkDREKvp6pUJ
3Atyaoe+ScrAka/GLwVCrrntFR4szvM1j3+/izZ7z9Xc4FlkygjWtRIzPrADDPwRmmZULT4x5ZFI
g1Oex2WzN95U6BtKwmjNGlOvUs8qIBtRhZ84hxw7JHpUK95ojS0q241uNtOaEyD9s1xj4o7fn6Is
mtKjW6KmkE/Tk2wMCw52U6jcurg/N3eTY8BP3RJ7c+0IT2TJ0zJH8cD9gqVv9b2Mbi7HjzEwHL1n
Yy1vD1yQaDHpI8GOytWrUWlPuuNu1XijPCcuwAu5jVCTNma1mYEQb5pYhZpjOnWRJoT5k79hVjCn
SrTJxrPv+IR2jiZqEFLVEADRUsnoiys1OeMwjqHrjWIJmdnGZKR+ToYEC6RBerTcXL2OacIO2/qU
UJj+8TO7vtnc0V2ByobKOU3Rwgh8jsyEcFRipv9jthYp8yeZniK8LKfHTqwVZ4pg91KhqOcqeEmf
5u5csc8yvS88Vux4Atdt16eVKF6p5A70wRFMNwMIDJjn89mdxijAmFqcWdD9pIfi8rofmoJHSgG6
7KyrogTFIbb70VAFhWzYksXMnmvDLjdBgMW9JUBkp+FspB0DoCIVl07WVUB0iN6oQQB3VDjfVnn4
+1j52/7OPwZ8zjB0eR7X2mD+B/JdbFIm5eMlsXdt5PH6W8GRnIIuTKzniMiKIpCdWSzww+owWQpN
UI+9IgsCMsBVeQ7avNuhg74ckKW4P4Axo6mDr6QjtqLrMRsAEMkeP6uED/PyD53SUvjDLIEbF5Vn
CsVfDyCDOesaVE7tjAti1A9lsI3kAc83qpzl6qswaznsANnKeeK0uG57/sScm6ayU1ca1kJ8vGRA
vIylfUKhqe0QtpP2NFbXMV2OVEXDMCHh278snK6yZTO4Yr/tFtxhiw7ZANm3nvlv5UXYiFUILJ6i
NcL63gwDznflM/SfEe7Fv1OraPH/+O8Yw+vVmkM4ssAVwQR+e2tAjv8tV5XiLP9ihyoMW65QGCxH
FAF4jOgFI/yad5qh1gkuIP6sKJECDqG8vgK0ioPe1kDjOE+uA3XcDRCzxoICDJexPfnEIr/R2sgZ
1FsJu3bBgy0pGi9SW/wlGQ9MV4evQpfDrkk36aQufdkT53GRnqqiam0WIPq0bdnUWgKPI5EQ00iT
XQgpWwxrVimfp6BtHL5JljWEXL9umN2mefE86Wu8q74Fe1+MV5fZl/AMzNdr+vtaKJCwlyw2d0p4
Kqtjr3agJ/6xAI+LjvEtZan+d4xP8fJ733dT+OlK6ylY/TGke+UngmlGNbpKWMzrIpku0ap2z7Hk
6mn5xY8xqn+eOrOA4EE7ZX47cQGkPwtAadMdblzlbnUvPoTFchqNqrcdgrhPjDocWUR/IURxSWdD
63cUeaNQ5cC3G1W901rYm5YvHITIp0bIRIDMwWZtL0/nU15L/c58ukjSWHw1ljLx0tfdZMsGlIh5
Bk+d8XpLexcw/aTlG6Oiqi3o7B2O7ty6t+phJxKaCkNikBHMfWCTKBMsPgz4ayCWs1t3yDvhfayK
76pfXORGmr7U454eN/VoHRASUTP/xJ/g8YXi/471JNxBl7QxOkaKybpqKMR32I4/Sy8JdScqWPRe
4jIZZ1NZ1hzfTrRiLDgpHkcr8iR31UutYTGRoRghMMH35YMdpaa3NEFQx7tCkuxRYjplFw7cEIL+
4eCSEumUFpM0kHwQuYCrnN0K62VTZL3TWbI806BWK66IfI6WUGkTy6B3BcjjUpc/GswTAE92UOnh
fnRatC2r9+ed6KyCRmWMDuZ4ikOWCx1ApgDg/J3hDn05oHWwKoIItsCOiO7q0nqUeZcARJeSJ5z+
PASlm0u9f+gr67KjeobsDzXuxu/KHSa68KDtlAnhDYl2qEpGCaxhtGEKxyzerZnhNB7B+XoUgxP6
k/3lcr2SMIQFp52OPWYuTLWse2p4wVaBgTdIB11l1N9EXYf+G93CIAVG+YykjYAjHoVv8+aAkEbS
pgju+YLRR4Edh3y0S8USz1A9sTyTHD6u6U4a6hkr3aiOkA90owwZknH7YbrSo7mW44z+C61hxm85
8SNnHHOcRs263vmuyiorIdzwVfyO35oJ3JbedoHunWvZD/RA4SnDb+oyxdWAnikwUqrCtFle2aP/
/VM03dgw6YnnfITeA/pNuS2MghIcGJHgJhq3Ts8P8rxlnjLJC9zIOICCthSAI/pm6h6GD03vtYdi
W6NAVToOyntWRi5kUCJ3QW5JArmOmSGroMhgucdlzFl1rC/iKeVXmRmO8M45lkKGUMQhKqaWPOQY
V4jmZI7BORDIwrMLmJYrop0xcD+ixsZKoAMNp04KvZl5p/2d1BQ/e1SEVJ5SsLfmrWyVbFijbUXO
pN/G/AhGQ4kVlq6OzNVLIanIsvW85GwYl+9NaSBfjyS+fCIwbbpohWLZnPoLh7t+z9AEH3TiZjzi
Jfloeu4cSI0gfEMecykyYB2jtLYd8LpfVOzH5Hpmgr6jWg6WGf/dAWONFXU0MMnc8ZFjejE5lV3e
qFevruLIkr3fWnyn+3qKVqcUpuBBi4WQrTrgy4gAV715QfnCINIfYstX4IVh/V2t4oGpxLpMPxvu
JB4xUdu33mvukFrxjmSCFGnct4aBDnjya1kjKBfWP4eLo1cn0w9ZTpa4wfXiawpr58FJSiLzmxX6
TtgerdjVCnspKGyQv8Z9twi/LLs+K8GX3aPS7p7EIVkrvbbTWMr3O6WZNocHhAPNDESjCygNMgf5
/cSudjxePHVD+TWlJXlwiO/pfL8wq6s2Zd61rxpJ69sBdxWlwEVhrNTV4SGCIXE4j7i28ZR/Mh/w
VQmAxq9QnJs6dEzCAQqjUGwq+AbD6tVn573o/tdxYhQe8AOJ7HjiZ2xRSrQ9HBDGBZt+8OYB2jCq
b/ergnYp4cItZBjT+YGUZ+4D79MYI9bD18Vq9TWvs93w3p3C2EFvNlRvxeXEW47y1e9hq1ZsGeZV
40pfPUeKQkwSP37IO9BB/tKFk3uDyylGTgdEK6dmtpzwbohPOaTIfMlC8J+GLNtZL+uMx/rf2tDp
nLCAeOvXNMPPYiDlwVXSuRb5+8nXVxwO3yIMJfevDNKiD28WYYgwhhNlQ2crPaJzHX14rMu7hEgp
76pQLwtpoQtH5caqpLbHpXHoIQL7Xqw6pVLX9MMua6bwc/95mQ1BXnC9eKI0y4s2Gr/5ZE9aKsQL
Wi/SVj+OYBPsd7P83a845MsFlrdugzb5gU1vF2FMpv11YO9V3G+8kVwr2uIHYcVl8z2GkE1N3r/Y
HzqXzT2cVwjFeK3xNvMbp9gjpQ26uoeWqU0wDxKBOWy6WUQCbxzeIF2zwtW/4tpCshQuhwB80mUD
4gkegSzRt2/XoDV68LThTrznxYZgcvO3tOGdCE8Pk8Wue3f33jxxt+g5E5YlJs99tzcdcrk/FdBi
37abkX/Y22kCzYfoqWNEpTxAHIyC2Ucn4gEPse2l2J4OgxohrMTaUtULHdEmXyLnWxvldxdmRXT+
gSKJDwMvKCeAmNUdlnZWlDsx3h70y+R5MwDrnFtgIIsM8q9yo/KJvxhPCX+6GrNlt2ASpTMAfDFB
lJlcrwEU1Brk6KihGnhaEA+djX1kuxWEbAniw5nh4Jcsq8KstjWClGe6RxSUkuSchoBYmqCQGBP9
0W3m/mSng/D8JjBdXILK4ESP3ZbqGqCbWQxx+20bdN+RN8YKO4ePIMHWtH9kscj/YDBXskrz/oeF
0qeVxibYnVldMIW8bT0o6wSO9qgmWUSo8vXKD1Wi0t6XQKIVjVz+lGDbHZhzvHfFt/v35Q0govOs
c91zZhInDk8HAEvEDh/77URW+YXaqmSwSEnq9ZZkQGfpwxmhmDqWCm5IKVXbr0UrCMMqM8JgELKJ
3aD7eKiFU486aef6COCK/86QJuBVsv5GWtffe5bY9J+fXpb4KXuz9TE33Spd8ZASIxupqYAL7xFr
2ugO5iD8YcVmdMT7Gwi89yHLw3TeNaWzqbM7RczXvIFs+2wW4PkRLeq2NznlLXfx2wRDN3wj1EKV
HSUKdDMZ1PQEQDEdtGoOdIn0beJnUV02AFRW8O5dgRe3OS8yxQ/GkcY/vZNIrBWxSNvK/oE093S2
t7OUqUdkTS8t8gtIYAlA693XY16hVvO2m5+iepxaRigF2um1VzD0sscIex0Goxia1pP6dwz7WQIr
R+rMLLSxZjeftZmGDm6lCjLwObauCbuLHhRq9oP9YdL4zQI5StGfhtkNTthdppDvGQMLpvcArlgQ
DU2wUMHQRGvadMjk9sj2r78HqwzyFqaSZIkia5JYlforCBBnjj87MClCW9PTNLGMKnk7aMGQJJCj
4VXcxkFfIvjCUm2jjz+Y5mvDm9DjEp2PbbD449d/6/CLt1oNbg13QMQccc4iwSIUdpXGtIt59Grx
ULfBwIplQ0GCg1+Q8vrrEVohGBvKWFUIkjEnl0nHyOrMN3lb+JE8o2rSqYKjSmkALiKPBhQb7piL
l/QSkIJy2UPtXrxrKKsnjadfY0bmCU35F9yBh5gT77geSMto8f9iiUCIiSRuKLZE0GlQ5DprDWS9
qQ9Yx+h542HCw7izGDdVwBSCtxA1AvzxL4dmmo2BnUEICukoa4PitkbPyCnHXvpI+jgqK6AgXSqA
ChWMEgMeqTtPqPi0A6XnXukaZrrKl0H6uh1Kd7qQQwhe928wHfrgt3AWytTHyxJMujjhumaUQKEL
lx8PKNm3a12dxIrzKDfFII4s20d1nJd9FU/Gy7H/TsZ4aNNA6HlwLU7A5DTPjZY6Dh2ewteYiXfd
4H8wKXj+jxbYPcRtrgeSwOuEOqog/sccWz3HY0MrhTi0KIywr8o2UMbL+PdM1xcArTjlTUUSsZNm
f7ZO4k2hqdpQdH3tX/OG04U3QIzqknTK7HAmTy95Elm/gwm/ByOx03RhYJ1qJCe+u4pu+oOrVfpm
IqrV5yyWsY9/okhFF5cbMlYBdAqrFD86wu/HL1Y7c/879P01GR8rg+VFSkQ4LAmyObtdjbgLMHNa
/ArUrV5GCj7MjKGt/dnZGA4srKeFfnKhqq5KTiKFWN1MXAhxZy/oUbOKtOXm2d1+C4tNginyflgo
dnRp4g+SoCk1+9x4CprQcdR0NmpXzr6gaIPLi/hF376jVaMFC6neo9+nZVjbVKGwWcbRmecDMXTf
CyJCXbzLSjt0Mecwp08xTSoJV7md47vegzLBjnCxpsnnJRcYanaPY+cozJPiubh73Al0fqqoyLdM
eLKB5T/NWq6pGl1PSUpo+SUBDHyxh6F9QITVZj9o2mRFwyFwvCMjwSufAg3oUxvWyoWIokZr2yZ+
LGBqVYi8Poe2J8/w3STEMi+9bF4lqd+T9IEA/thr9swdi56h9/yzQVauDcVOCVX/zZpzawDt1gJf
nv5eB+QnpGQWvKq5hvFX1iQEQ2YW682DYifhtEVgxppUgjiUuPuGKZak4jaxaHCHNdkTmCtKVvq4
qn+9Gv88I1MCeT8hzzFeBC6B3Um6Q77Wr6OYtlq9VUPc9c3ecBH0rBwLJdJ73yB6DCF7BgpL3oWC
qsykY1jaJc6fjSvGZ6gzPTgP06IVQr29nCvUNv3M27LkIxvVd/7/45pggA7eoO0lvDuZufiY398O
DAzrNCyyeshDJeBs9cwM9i1vTyJ/kYPWyz5vh6aZs5iotEgqgc2T3rykZwvBHYZ7L08p169nAIkP
2P75XPnPmqYx9NRuKZvTvynPKpxGTfea9UQHl+F3BM5EkzaICs72V6bbRVppt3bS6a8CHW8gN87j
IuyaN1yMhnz0Ux8M6WPotR8bgK5TzQCrW9zi0vtYxO/ymLY8qs7WqnClBoSMSZ1qvHYOgplOY9gt
/qXoZmvMqvo56uw/TR2wtVfmmwRkZw8dxIH6IyLQ8rnWMvpgGt2xIehMHLucdywuFEtQWLhVHZz6
qqOPGVJGpItMFw0sH/Ty2IDFRmkNXmfmYqxUz19+c5l4fSKKkfUuP8C4emIZB0mv2DfQmbe4bcKh
/4SN3+c2JvMrLAdLVlzwYyC3jzCMq6GApJLUkrObyMFe4vwtXM/IKfUoCiiPJWtzOi2zU1RoHU8a
tnPE1NN8T8QLhToJvqZ4uU9HGynEn6a31NX/JLhv8WRyrWfdF8R46O4KyP4DRPxjHCz3T35je1o7
87biV5PfPFIesbMm1RgGJfSE8YetnQOQpTO6TvYsWjndwIJSMtdOrhwb4LPhTMbjlkXUbyIjc1vL
sRuzwRbkVGKmDKbQcDUr9746foaxoKoLRY+PF8QG6TNeAaCFhKiBVsgQ4YNR2S6KwIRMYrvT8J/G
0+gpnfr4JCRGCf3wVvmDQp0VxjNPQazzXjwxQo0CIzLUQaLQ53vDu6JqYyrIrTFEHwzFiyVdZojX
cJDPYZiodRbg3YUsVvGnFQBR8l9pXFO6Vf6NAxfdj1wlC2dGmEjlGYg5dxd0qN4bBv+WcSX+rvpQ
Buts5rbYxUmZTCtv8CjfIBr35XDLAzPsfkuLvlTbXxkBhq17fHdFLa/B1InMwfYZVoT+4gmzGsFy
Qlt4YNyJ2RUu4L/b7Trb9GPKRj9+UmJFwWLMpL9VSAaJUoops4s7Oo2lSUmfjFIZTDMalUIYOcb8
4CRBtGPyMx5lHfqxd072T3x8OHbqrX+S/NhGNcvd8B3OjGiIEpcpTjWdfciTqk1o+NTCQr+NbDhX
5VLiWh7vJcXaQubevKs/abXe3OWGwubIzHUCkBhg7e6B5h6bFqEvbw/EfMBdsur0FCUbgidxm8wD
64OzBxM+MecNI/eAVCpfztmilS2oviRyaNNspo8XcuM6fIlKLi0PY5kc5WSbgx30h50AbiSIVKIH
8s21kaHQP3BjFukARPsUiGrnIbwWhnSTccn7oJ+7qMkcDyXEquOZTLSUEeSQzqF0klKbK2RPJOGG
LiUr7cm0oiGkC1GkR74aVdFPM7oSSUs4qRqU3vt8ViGEutlNPzOUn8AzTs3YdWJ9TLM/jquQsweb
AJO7sT+KA/4rnt+wFdqsrH/TaCtfTCjXi25dPj3UiPpbB0v14EbXxzz3HO5Dc283mKhYYOTjRXOp
oDkiUoW3UcNa/4CwwrZ2fh+W8fCGzvWwJorYWmeU8BAnnAvXx5muIFMw0CRHePlBxHuom7NuVFt9
cw+BilXorC+enzO8Wo7pe2DvoslQQs7kH8qLDBRWO4Taor118IX8RTZ25DGB1hpvChrFcMDPQn5K
6vGg0VVZeL+oTs6lloIfnwYs++QsFJOGubgNKD7nS95/VO2q1xpfSl9yyf7jkJrkVra5sUl0om2O
I4Th7CMPF5a2OBimAY1kUyQqW4IFMZqvkmwgA3e6g+FEFdYhqNZ/ZRMxqfjL/jZAXB3MB7F4Z18w
d5j+5LqfB3lx8KulsmQH3u2NEmDXcxMyaA1bxU3DEOvTjGsIF1psF7rw0eQ5cBBAZAihDsRxqDxE
ukGTXpXHeZknT7asKOJB3aHC4zdVSuuuP9Js8RLtBqb1Vg6WKuBiwVkHfIwkyozKJAwPNgDRFIpc
CIYcR15BFbknFU+HaRVw0qg37Z7COAHN9WhzOUulrc1HhLvX9yc2sLWA+KI0jq2+Aw8Q/SyXanQh
numlD6Zial5vo9ntl7hc+r8mqAw8pczbFDovWh/ICD8ZV83E6mpddMfrsTZa6utKDZjpgfYHeUcN
9ELmfcw5p/b7wtj8/pb/wl5GpGgkllyMgdcXvcmuMWnXtAdsr8V63LDvbCJ+OBsQPEbs0/xpVfiW
3b46n9K50wFXoQtJWJrmXQi20qghX9ONnI8t6+xq0rIxUJ+WDx4RK5+EmYIjVMh5a5ADdCOrinGA
BATe7HJI7aAuAJqYBz734kK5fEmb+7aIYkJHCcodJZG1wLkB8TS0dww9s+vz8+3kDCWcG6zhqLa+
CAIH9F1zIENkP6B6OS1FdJ95Q0+HpJyVilqf7SAVarXFXzNgDadIyRjXwc+xEYzBQxcSpIOs+D2G
q9nNSDcESozEQOTBM54E6gfPNyTC2fudx+++kDJMoUtBvgVstewB5diM68+5ol4BHwb1CRwQoxzY
xJbv+po/RpJS71bk3JpfG6VlnUxNPBfo+0j5kpr0NYoYEgLZTq/ZnhGOg3Wq/JGnDRCmx9naU+Qr
+8pFhdLkwmNmj1PxHcb2htM5tGTJkbg9pAHj9vm5YkkR+ihFaDqKWeKEEgzlkhvpGwuQ5R6vZYNv
zi0WIbpaQnE+YNWNvS7R0RA0ScAEDnOPJMydE8/43QYbiaftwjwlFzDsVIT9NLbGTL2JyBhcuUGn
PgFS6NaItq0/EUVbXnoV2jHiFL2R7A/E6ZXZ2clDP8HESH8PZ6WRRYJaLezDog3Da/xWVh6ev4PV
eUOA0iMLdHhrFJwgAYtR0vz3XYqiFaJAKOyPjP0YnBxxp1zZ2rdqaH3quh6HJumrNsyYiUVuU3YH
vZdi/ou6D2lBVWyQ3L4Y7MIfa6ABGWUS0rShIvV+rnA1FyYzLQhOD6ufAGAh8i6YlnyTkE1m69Ei
8t9c7TFKoI9BF6Jiil14wNFPJHxmFRd26wthOlfe3UKBtAUmRS46kzu7sJkzO0CGDC/6eu1g4B3d
52D44c2dsH52A0SZhCjC0sb0/q/5f4wf75qOiUpCijWTcYRgOa+kArDY8Px5GBZPUPzInDawC6iv
gT3BjwGdEt7D3VizkcreycyaxJ9Cjf/Gwboxd8KXA+PeTYRBGNWszZbK1AV4CvIWlTQ/B14WOBc/
YfRlyW6xOdjhSR5YiUhCZFfNxG6YF0obQVGf3OQqKsIMS31iCOaLuk2b/88nEiaBP4N6xnQuUKhO
2x9+iuVmqLXYcnsQJF3JmIeTpifJFCPjxcUcGoc5jcWmDEmUmx8bmJIcqmchMxXl1zkq5tXJktA1
6L0d3JfBejTLFCxyW8qXwqcCcUxImwt8UaOBty9D4MucvnP/hL5Ta8Bji1dpnBt5raX43cu8mefJ
/W/h0D9hLPFx5st+DfKKXyxMxz97QFPZa5Gjhs/nbv+R2NMskh/RBLa/dc5RktMG3CIryQyhCcMm
iOG96nAQIL1EYQcqQNEfiNkGCJdCCveS6WUiu9EDqN+KlYvjF7rBCkQYhd1Y6WeuYSC5UNaoRDUU
mfXCXE9U36HnshDCAzfkkhsLp2R+oesT23auiFQSfyjUNE0hxjqreNrHOPSKzwKRN7OX58rIMwOO
cFDXCKBHVfEmrQHU0Kj7ZXBzpVT5SdzHnxhXTY9Lr1hiso0HBbGpakMFRVY2hAWa9b2tjvgld3P4
/WDACJSQ8xSGMVm8toleq5/WaR+e/3kAabZHjQ5HSo2d/gxKX9u4vUE2RS4e5/Pkkccm3BLqZ//U
bJy5mw3OAscjVlDmRCiy3WSG/r4Derkpa8OTnJXyzVRR2G9gm6nBoP6mFDYoFR53KLWcpXg5Wg4J
GrU6bFGLXxvaB94Y/td7mo/TA5auS9ZPnpY28A7T75qI70/9DBvNrKxSpklNW5A+pxg4raqc+COi
07PtVnCEEfmUd/LIIpTruyeIICs9rYvTbMffK40WalN2Qeokp2qTyELA8/B27nrE2WW0qqzcw4qj
/DQLARqrPwdEmdK88W8FxBIHG0i7GR+xP5hlXTHv2CT0xDio/Z2aGU47NyqhdtZvIwzokbGXAOm1
IJviDVTGHfPpjOSXSSjhRBx8jg20cRhG2kva09LqtjGPbOopdUVjpivsm1Xi4ezUWHBt5QVCCEWy
dYKZ7ci5XeFvhWhnF6OTR4QeN8xkU7nyB33JOvQpo5KkWoIaGmjLPA6T7o06oF1PyM7ksiW2Vr+b
n73iut6XAKfuN6ldhQX/jQTqRqMzzOBMLUQcfyWZ3Py/x6MzHbbq+eYk2opF5B5AkvZI7P9c+AEW
00syFHynGKQh8xsYNTg7G+/hFUPnw+6AUwXQGZ2Ko4xYeMS3Dg9M51oSoe3Zm6VLDzxZwcXgJ6yv
6+iQttSGiRpf2c21Uf7HfYu+g3vhtzwNyUUODv/wzu3uzXTU3ok8JnfHm0Q7fu1e/Ps7HIwE43KI
j9vGvO2mi+nQu8MG3R7dNHxI+HiK7DBihUkS41Sln1QZUP+g/9r7ZKQ/eL9J1vmCyvZXFl/0h7n8
rnyXQ0Cy0m3FJOrjXPBngJL4QP9hwsPXQDn2fSXZw+cgD0r4C1v78SKSl8SgyyTnlfaL8nBM/5Bi
BgvC/GOCscX6pc+JKXPbc348xp9GBbPM0jgKwip/MZBEAsXht0UBNgglu3/Pi7DyvI1QSb9QyYhT
uojOqa4egsUbfyUHjpXClLoO6ynXm++SMbWVJkV3F0DTvnLlf8dmF2iXeqxH7z9bn0Fj34HnJom3
x2vApETEBzXRCGfGnSp5NnfXGV+o2QWwhrmGcuroTXsy54iU5gfUmBf/gUFUeG2aM7i0/GD8tPrP
Gmq2O03snIUWlI+Yu2olGnxgFYsRTmoeMvQ2B0LOOBTwL+eKPY249UjfTK63wP30ismpuE8cqd6X
puIcrRSC6nzhmbR+QEuMS8Vdfv7nFNHqB0MGXmJSCZaXhNjFVK2Q3XheT8myCFNCVFLseY8t44WI
gXlxmbSTHN+J5HMOFzUlHPiehKFw6251Movnz5qE5rTIbGLNxLs/CRTvehogNzF1uaEEhsinTGLQ
YMm9cazVSsI+dX/3ri7Btb64g5r5kr61HzIgElPyeiCuAphFGULxEVxUSff+L/8WrfnRy/g+of7H
6KMbsu3WQJUEwU87UgmdF7hcKX8SLp5bYUnPMRPlAhGjgTwOUApKkTvl4ybFQLMyPn0t0ZkK6kvm
OMhvEB4Gwj/PlNXKAkkPzQfd/Bsaq8hDfY1M5ZhHvNDkXkRbGR3EHhUB4kJPmnqw0UZBxdR3wXQf
GuyGKqpnCcDwCDNWRkqTPgJP7zNHYqFzzpiDpMMyelfG77QL6P3JGSAkObcXoASh0OgIO8vV4nFV
otix7diz6azFlwYP/A9EhaY9Qpf/ET2L8K7++TIYBOoGqbIISotVAdKQUbBek43cInqGIPqiImJ6
NWMw+7NHGMEobbh+7TpRcAUg3nWjtpQkmRda79UiEdDLA6qi3my9VMVvQO/wyhMMHmX2U+8ikuDs
8nd1tCJMFLGSgg1FqnJAYyqIpDCcyrEwPCT8/l8PPqtDVwCiq5CSGX9CgOBOzEn6YvLk1V7LYeGf
hV5FkWzjtQek7j/y/buPPSeKDYH2HbmO6VPeJalTWr2ZgPM9VjQg1MCSGnB6mI+9OQoxkUfv6YEZ
xBCHME67FV/bL4m3z60IIVbhs8Tc0HOOQ+eYqJjwcXGB8v4M1+5i0tejIWtCZxbiVFA0x213ylJc
dB9RqOugkW+S445jBTuHxV8sqPyl5h9fMcwTEC0vI8QJzobUbU4FidgbcYT+K9WSJ2wUZjJALu6F
1XC/gCVlrfuOlsaixSk9pBfEuGqPTkiYKT5hPjSrIqyeJ2kr8e3y0HLe0Uw69GQtr7KrNksAb9VO
JAnnPy8J3fjk2B1pMoj3p2SA4QlkHr0oAPXc7R9XDDCbvDWTGTewpRJkuGTgtYb8JutoyzJlzVsM
xTm7FqCusuhs742POeDV87MRRA3/cUDuKzUv/ZBaW/7mTuXrDIwxIWKNJnkvpRqBuO7/oHSN6ww5
ZgYPzwzfHyU+/6WVRRNZrH00E86gObVwktvtu0yfRCUVfn5l/Z+TJZklVkTKQjyW5jp5Rq+sBWmq
zZgO+T6qT+z5kr2z6bM74RKz99GmnY6Q7xePooD1l6q6oVsARzLtJ155vUGKcnRAVswJyAovI9KL
hfZ5sMl2V1T6+ffyZf9FpfsLxij++RF1zr1f+0WREOpluJcVK3qOMBy5b3V9ydv4Oqp2tC8/mjPv
WubWmSn93qL3ECOkExg2mvYI4+TwtaFuVUqw9FEGS5lFtQNCEpUCNhW/6U15EepV030imJ6yu85y
TGvNg28lo3auYSHR3p3OBEHY43CRYGqddYZ6Tv+lqpG+HLd1Tkp7bH9Uj1IL5YUoy3rBAK32QFwm
zsng7e1smd9Q44vLDj0H4ccWc0vkMi+4rCz/6suupfTWNMm29/wF7nLmLEqdMTSdfj4HWxXCswzv
ytwnS86hZhU0F5pmHY0lNC4ZePKC+Z0Dz89qNQKMmEpFTxEMvys+SC63cGvC6+8rtfPA0dyUmQK7
qmaAXSZaNc3nr2HD3eN6T3rourIif1oDnfbJWoLn36KhOUVMHmxrB52+aj66DJx4wEOeVA+sNGjr
r2axn+qlrn7hP6tLO+o2fPJ55W28EuhmPBowKpKDNOy+ZnDa4YB1bwNexFWAKfLbmAMZB86/ImwR
53pv6+XJAUYR4ixCz0smLqPIUzg4NwKfIG0hhdxoun6cWa12vAJQio/pSuv/cWmcsHWcURdM3aPA
IHp/HNWLve8Zk8d7dC1JJdqGarmYEE0tWxQEImQoFfgqmxCE161dDbiwXF+hy2NYV2jBvnhMfV7R
u/P9S0iie5ssTSZmYyWhc3Tt7nhdBFyrMzX+zo3nkRV7jr8SSc37TKUSkoh3ZVDThZ6w2WrpRh/S
yqi6CAKIVX3Nxct0hslkIUEKwLener56fDuGu7LgCnUe0eBhFfGUCwH2A+RHFXoHT3l3F1U5g4xU
ihBtcysUO6GRuiqMmAeb4fG1D4fXP3nW/q/VZg/xNlYOt5WNCqtiVqGRushXjupa7MIBsc3k9Z5q
iuEh0dI2nOYIMFv2m+sFE65I2q9DcapRf24SzKwv3scsi18XrCdUIvNXRZTf9+Tt9a9PgUlJwLO+
EeW2DVp+j9Tp7+IWh/yU170FpZfrqAGPnage3/NgCJpJVA1qAVSzdF1H7abgq/v8LU9SSqPYtGR6
EeyjePsMDt7ZmJH3xhThOACQ9eNRAIBayimwR9jrnbcjf41S/DQuePpHnYloK+8eiCes+Rh3EwQh
ntQ4qkk2JN+77CjIm2UrLnLxcx8RGLP1XbSj4mVlkHhxDRRuY3oEma5jib5f7SjivXTtTY4tOw10
16Pg1oyCIAHqCERbW2nmxmy27Lj81Hs+g6EjzFVdt9cqjeyvI+r1SntdgamzehvCq5+5pBKrKoSp
ZSmafzhXKfVzepYUDcV8jOq+fBwx8NPLVi0AthfKXz1HAw4BjTULptvbRHkbb5XAAaD8SknHku2k
wpzTSdTArVDtBoDqxs8kvbYAb8D/iv6XcrB2uHT8Bs+aACQqNfeq+8+mjyfdYqrAuG/dVe8qKi6H
nvzb5aowT3Q19qw17u9ix8ZEUVxOeL8Zz+35CmieaxaeTYky2vvvZzmVgoqUhWZCx3hD1lKr3Jvn
rgZokQq01WtAuD+S3k+OOUL55CgyfHtRNXPNY3biIHwpt7LG61LEMqlMfnZLKEOTdzRd4dkZAJ3p
Fbl1lRmhJNQ2cH502Mp96cjfNL+pCb9FIqybRUduhiOCzLmTIUPASNl80s1uxEF9yYeIlczbVN5w
Ks9RMnBa0bek5Y5rzr4Mq5OyAjRAItqXQVzLke8KWriuh5wxWjA1PtTMJjRuaiatlzwjpiSIcQjD
BrzuABHhQDoGQu53/c3Y8UbLW6OSvLzJcQKDGoiLEG90vL2CU/r3Xz3riDZMs8bVCu/e6rLogRWe
ip/rl0MkfJr8KohhsAPH97RFIaijCt+JYgiYmZiuMp04I1FZLP0/yOR3L0wzLiHhZNIhErbFNkuU
e2qXpuDiyVhusHgq36hL9ZiRWF8gF16o61D2yv4iXCR2TbLRXer072jXTJvtgWhYkzX3ioNjQi7C
V/PhOYHEQ9hgmAX5d8GPoSbwLN+LpLOGthSTmXErgSZUuvh/DMa0c1t6AEuCneBr8nX4ZYPtNGvj
EqQ8yixsfOeT1cazmYodktmb1Z7+ffXqjgIOj2INdbQeMfVMQxlAAG6cWE4y1yJUgOEIAeMwnXhx
yK/XJEcsCeQ9l2Ty+nrrRuu/L3pBwZztbvnOZ1j5wG1g+o7nF+gpA9uHp8Sa8J+twDcIk9yupW6z
NaWX0oAL93aGbNzSzdSQxAZp/3l1vfKXM1Dm4iXE6r6Xs97qZOWOMMXZ/FJ6P2EQlcIArBY6F4S+
nwI5BYNL1Zf/0Wa4J8MywbTDvBmmNPDMP3WcdcSmN/Cv3y9rqHd+DktodC4/lShE3cxD3Zccq6eg
nf3oMKJyfgqbt1eRHx9NOJxHiIHRQ1fbRnvgfdnQ22A0fUJrJ1puMXtzj+tkZH4v5t5Cz41V6NJU
RulN8hBCmerYeexFOOZ1OHbs/0UvU2OVKz1nIzJ0QhEl3A5ZvSkPe/CeuJMrzsqAl7Suvqlxir6t
Lj0jZFQHfIgirHgKJm+zQJr+CNY4Xk1T0RgkGamoiqt40xjGeScmBvYFmAmlX7d3fnHRUPhQI1ip
vTMG8fw85r/EJu7TKCOlzgXQ+xNBdABZm+Kad6awI4Gxm7kFL3NETjK8myPxeirnZ51S/dfmOJbQ
EnYYu8rgBcNs15RIIFyK2a6QP4OJCleHhqOgzJ7FPRKk4JTuoTPpkn7EixULidFDNPuGE+dYbNan
l+ekKRJrNWPled1aOni4reo2ozEs3tP2GHnOswdHGkyaaUi0Dh/rSyuBuERAXqRfm8vn4zbyHu24
7G6IbM6buhE86Jk59e99R79j2+UEUpF86DWvfNPbZFuSI1THFmw1wk+ERvevyxxGwpmpHUeklxQG
UeB88XhT7UPzEDHUnj4LG01QbyDu/mSbbTPJybr126jNLKPhbhRiyuuKq/7yYDXIJCB1gtFZMJr8
uFYLQIlgp8SCXE0fyGdQ8fzw3CmQPMuazhZieoi4rJ8w1ZTRyzJLvd5ryysRlSVph4Imp/y/oauj
+DEFrkMBUsf3sC/bzqfw2o5zUyFZ7ptG0Nw59cVk/dczMtp/VaGqz8b+ffk1hAyaHkTiRZLnLCKj
BqDQl/3oUsrdVO6kw5cpLdCQmJ6Md9RGQQ4FOerKV950ly3OezhkstnNCsv1ZCcFEzPOLgUabe/W
IfKkcU7gu4WA03JHzs2RVs6SIDI31bUCId/ct+2h2bDIPDSwlma2ydIoYQMIgWn9ZwbuYfpknfH1
X5+JKlx4PfwjhrASAMxi33ew5Mc33gqtddt/mUYwG2PRuRz6oDainmZBXzbwV3bkFzAhUe3UhrU3
h0HFQTzkf2dp2JxMrw+UYA/Y3FlRPb7AB3X90hou03NzJgc6v5FUVCuRBk21yGCGIGLldUEPeK9F
1e8uQLTL/a6bf0Fmll3U4lDPjwocw5g5lzCeyTmyL81szBJSbSFRiH9gy4OFdUX8+ocHNimJfE5R
9XbuqPNEdbL+arLcCOYYZsxxbnn+AjLjHDwQ8fSdxuGtXkWGRMRIsDNSOT5x58Vn5sxiHccBghrh
GhYYOOZ9+6OJ9YHYCQxQ1unYcZ2xxCW0AAguyFCWSLd2NjoX3GMF+6YH82YsPUkaU50gV/hLNlPB
wrc3prsq0v1Cvvztvkug/fSTYH3JPCHEeeGUq2IBd7BFPqbpwZzwZQ1sTbbk+S77Uk1Hms5jS/eS
HwJqd16hYREbvnZVufEwE/RqqcVxUwJ/EUL5d1jlUFkHGRUsxZKofj30tu/U2m5Xt/kXLaR/0sg4
tqZLDlIol6s6Fw6nj2agLHB/YU4r7CnlYLTRKskueSEmJDy3fKFcjjth43Ruv2bcJrRFn0+OJcRE
pnt4CQMvoPQcVL3nvBhu2vkZRYGE2Po0+7pWNWXaRGwcXEQ/s6k1mpkCrE4P/Qki4+1op9N1z7Nj
P4qfO2qiXDc7LVPfN6j2gYR3eKV8oAEwT/Fl071yrApofi8zrfPh7/rEFdKHCnlYrNOKrE7SYu4q
XPrd9l193bqfAenOE7Kq6b7iYM+HEesZCVQaKagioY4JWzzd3z+aH10JIVNSe/KilygVlyqJ3CGG
Bxj4FmDl3fm8/9pnREI+HpmLlxyKBi3r44BYJmYHfFNJ+iJAtW73plkBmsDXb21j8Hr2sZfOUwrN
eqgJnKmILMYTbG18SzSiwsjuPB8u4VAZeWo9LiTASMHQAhRX4ZHii6PY0TjSJ9SYoV6y01R+Rsd4
zKXyqOy3N1/Y0ND+MD8l44/ErxmF4SgC/H/5qaKNAiLvKlHzy3uxirBXyNBw7fYVDXWYCiy9SbHN
8tv4Zwo0jxLNovxYI8yvh466znlf8TlbnE3aEA+uZ2VZb0MQXIICV20ts9Ska08G7/iCPYk/uZdn
5Y86ZcNLu0rXbb27TkMrxcYcb5yyTVPBbwcakWrHx9Q3i2OiChV6d3Umvk3Ydkf/nTBRQ41RXTPD
E/BqP+Fwxy36SCQm2s0IFB2pipbZ9kTLqBszkyL/qNX+PA+GJT1eZjnx+dTqM3+jtaKg5lZT/cA/
N4tcPwAsifF6pArfZEOwUbmyXrmmPdLQS0hOxs3U+v/tqMj+040wipc95o/LJwPANyrRhWv5wHl+
H1EqavjbS3Vcy59lLXuHf4HBi1V6fXIjM9a8MUReyaMshEVQmAakkl5VbjwsOzKrnSicmlfaLbBd
CY6q2G7hvQh7ZlLE7QXxx0dRghjvZ/iPg1pja2DDxN0SxxuMouiBNj2w8V4ogGb90hVbxGvX4yGh
rj16OhivLr5LNN0ExZyRKh3pkaq9VbLjX+mHzpm5DkQqfNeK3FHXfYXGNczTTszYdoi/H0cc+Heo
bcB2G/DfFotOTQk/iGVdzRi2GeFgd/PKEH80+z88lpQjK949GFM8cAIDLKrWPm38O0N96n4VCgl5
sAWwL8P07L7rCPNvbs9O45RO1T4MC5ygmX8YxZhnj3mvZYwwYUKydlvHf9DBVJb1Br3n4ZrfgGFb
LSZewt4j/VRDbjYWbCfMzuBWF89MO0y9t5q9yf+SnAcU8IGsjGb2juOPUBfsyTnJl3jh+V5bVsF+
cbUitX5Z1LHofMiNmsG6Ma5LJV92HcqM0K7BLUw0zsc/YLEONxoKJoSq7PhTKvRAP4JuD3Eo2DLc
5RSvxjLZ3BIkSaFnplJCv6Khho9eHAjAdtqGRyiN9ECOjhMIl7tnejQTAfnrItQwqBQy5CaMhlCG
AKDttq+oN9fCj3GPlNdpCFkS8kJRPr9LyHTwTjzgen0x9OeAzxXDAi4+YKg0dM9LaetV64yCnw7j
lboXJfb0arf3W0FwzDb62jlxC3LBA7OIU1en8lXtY0onEiAR3ujg+2FAYS0TUTokKKcWvHu8F1G/
1ybHIqcBtY3nZZpuzQ46iJEmM0LzF0SzMCaDbM0u14YN7DMngonjBmmfhuHnkSnxnNK1m/tO4ILI
UPVocawR1naX6eBPFtByM18UY5SItWPhKEj7BKmXnJjx8PCvAkg8En/e5P1lIEFPBjue7v4/JOM2
5GJXR87c6N8GqGBAZ4yhpF3S9UbYJyBnztQaB0Ui3hS+T3z97JFEDWKSquxJFh4iSw6k8auQTzXC
3Y7UVtXRCbx8tS7JnE9/zgbBWJ6ZghLjn+BN2iuUSnhiObauolovCMvyXlapNwZ892U8vzCrw/TS
XCF3Z3GGAniVfuOdRyO9WjNvI2TfW1K/wFwrljXd5YXtAMo2by3uIFcr/Fry7UhzNkgpyW0qAXuJ
rb2HcPBVUTjtCGZKqDBIkYVQaBwT0wE215qudFBDTa9Us+/XR8XDArRQcnQ8HDP4dv+nFMILuERt
CZv3OjCjWaznGvijQDDE48CZ/I/cb22aev5knx2mhy3BAgBRHqkAqD2Qq6KlLb6OEwqPpvm7qNl3
TQgZrVzl4FwV98fiIb5PLZkdaUP7JzzUCTMFU2RqVuPKnaP4rzmZEGcTUbkcFpJBmVefipgjx4jJ
MOHuayxK27tPOdTVcboGE53krbNAf+wq3gHwb+L0J4Obz71fgyKfiD9bJR3jSNGRTTngCquKlvM7
pwqAJNVrcMxiOI/j7eEfZ4VsNfMUITB8NqwO1SzQWwpN/kjwcidMGwhiOaW3a2gFLCfCNk7v2r+W
IqmacCC27uj5rGHhT9t6Nm2RHoFny/gdV3da/Gdjx1BxMJdWof1QpE3r7bATLy6JLEUzgyOsFBGK
6EVMUAQu3Fa/bwpx2utHYKAARahJeQzuNQqULP3W/IJDONvyn9dUju7bMST9jmXXx3K3nIkVVO2W
DjUBGhWvH2djnfblDCk0pfA61gKyoHCoS1bwG0cRmGTr12A+M5ZEEnNpwTrfHIZl8M1a5XeHQYsV
DVDazD3m+You1ELPj7QgOBjZKGsGCiwNPD26LeRUbSUE5B6RjXNNVlEQhhPKxgqXHi3CrAWn9aB6
XMpfwtx7y2g6ZfONRSt6fpU8UconM0JkmE2PhCoYWWhH+CZToeczxdRV2TZAsygx03AQyio0JNcQ
BFqY0wrY/xbKumVtvkw3OSlMxQfUaEqxR7U6T0/Ohqbl3qLREypoJNa68d17aYibUva0Cczku5+u
TZFueI8PJ/izh/yx1ED8zgMRYTIMGn5qVfUUprSeWh2edkqt8hSnPE5ZejuGmkvJCivQ84PEwJ+j
eqamGf2uNJKpMuU9xvhpmDxBaBNi5sKOQcCOuD1h96ONFRVmTnufP68AOyOy3vhebpjsZexNLRoA
ConWfaKtRn97XdmBb910lBXVaUlmHVNVCDWoj5ZmvvHp3GCa/o/furQ9LOb4PD6Gn7DjcczmKkdy
52YQ1iEs9ZSkjCqnxHj7THaNfFDFxT57GvcTXFe6KTPQuC94+DSS9US2GWzOJjmRKVWO0Pmwvqve
WKzuZRVqF/UDympfbpWqcDQESAm8kZoowcJoZ0O8LGqm2avUHFd+/rwd9PAzAvjxFeWoD1pGjq9A
fnWzu2ToepLmqv+fr/YsJjMTUwfD+/580L30jeTAtS0szR5+5f1Rb+rBb8oLZ7iRsRkt5VjlYJrv
X9qzt6NmeX0eviLP3pkOFiPit3PJUHJme+sxGG1nK24yMuzgjd6r5gytaBzgfT4umMj7XzGZ0UOu
2aR75CpVsxt0IGWr9PEDfgq1Fx0rrlLeHpFsyW2cKABncYsk6urAH1t2BpzQiLFHGw54qjHVobde
r9PvhkLBfjozdwo8dkC8YB3M9IhmWXAgUy2ztAjDER5NSV9aPwZoriV8HW65lV1xXAQNLCjZTL/P
T6slKcXCUjULMFG28dsVGfEQg43rJ1N7dP41EwrrF9bB3d6EWGSlrit1JDjdzFM8/4zQ9RZk9wK9
9tOzYpCPmzojz8W1HTbCnDbc1v2UmCdmTG72KVYucHAnl9Ps0fWOu5FNwlzbOwKnnxNyKMMPTfIH
Kg+KLDdzyLiK0o3u6C+g3qoYDaRvoCH+DhESt+kOCb1WAAdRTcmtEvuTHP2DlIVcfWNzpZSUNQLX
ZG+mzW+OpKI4TQTYGUJUWyf+VLU+Ut1uMKI1eeRlaKgWrInbIYVIA1UqqM470S/bFAdcb4o5cqT1
rLX6O7PYlqs3LjzjaIneXPr8np0GyPeIMrgpRM9Ckmt2fKPsmkjenDVFcRNTpLoG463h2tLOpfWx
6Y7fG4+pUtODfPNguCvoDIp71MPpllp4n/xx++SU0EgrgKgaJzXgCwlgqH9zNzFi6DMFrQnqw+rP
KWOUO/dalezANdrjmw1Sxd6rkBTxzN2E/u75GiOpRQIrC6bMbi47e2G/G1DI8F/ORI5gh/9+WoyG
KKVj2oJpViHR4PlAbMcJhHhn/rwrYIRnflr4/ueNrskJCmMynKnfoxMTqs4lCzKxmjsWloc3oREH
ovnX1046/qeibH2w6ZdCv6NbIAQ0V4fxvd+/z9+steSlEyvMYtgPJdFAeTox3Yp1kbYJ7CEtBrjU
RpKbWToiWAgTu10Q9n+mPSUua4HczWLTBB6EAX88mC58z2VOcU03Hsy5Mr68xCyTaBX72FrjPU2W
EJKfI9Fbgxcb9nE8LaAXwAJ3FL2/yjirVHrE7KkDuIzjZ+jgjvHxf3vYf2HhnTRBGX7YQw9r2JZj
lY52XMhhqx1pMhgUSTJIRwFJfwyCmrvH5bkjhCI/WUGglvM8LTfQ3Tc+WhxOePH5gSsMfhy6Wqh1
wZwTwy1DLAzkkjiSFz1MxSJxuzb4Tg96WEZ8N/aksYzAEjKVehkkeMxgDHF3uje5nkcC6feJXq7G
hc6c/n+vFxoUuTJEIKrISmL6NPIM9pVMViAmjFkTITFvChqxDh36T23wU/nrOOM8TtjFCkk6JQb/
hg3Kd2on4Q/6VNoa9gzX9/Nbglr+KZQRysguNdU8lMPY9fo92R+pyXXC+IwtcK9ooPkp92qzZxIp
iDJZboniJd2n549AaMk9PCTlrVvmgKLkmSkTkcqB6/yyHaFdA8YceCzOVlZknULyA9yCSm93i+0v
ypaeUst8osQyCbbpD65C62b6E0zqfmyYtVAwMpjwniojLvsGJ188kf+HQKN+W1iQYoUea4Qj1du+
4V9FDlRDX6JzogOaIGYKQ/2SaB4xJOF1Dt+95UEEMN/inqyiEpX7MEbXpMb9fsgkzfYp3VIeKzNK
lElFfYmUkAX8VmjTbe2YRI2dkrHXWvNd2T8bua6XwI8br9sqfaa3pJfwsD6+qgVstlGnZaRAnBDH
xfp03ZGyQ+rtmxt4BcLEFSyGXU9HDXg13IG3GkC3Cmh0iCmmR3R62nBdVUrrk5bX7JLG0pVZPP2y
ZfaxfpBjzWFaeYrLNjmVeh0Itfm549n87FbAa1sgrlSlx4L5zL+SBXZVTG8gxkiJ9dSyFL0IN5uh
rQ67AXeTC/SsZOPWJ3ZvfM+cOgqGBvY0NGjkLpYRIgEb4McwhLSimM7cEkS1yqo38w/YbQBeK9MF
8QbxpwZHGKH5Dyqx7RskCXnasyZu2irjPVvJeVgAcT1WvVehFx914ZhOslkt7n0MPRcQ3m2dB8r9
6ZYozlAaAqiwqfMS9h4HxQYianQOE6z0IHENwXkz9lKjqAb73AU7IgXAvDhun5OpQPdVYVJ8QWx/
akTELTBsNexfAHcXXN/DxHoEEISLmQyY7yndde7a/TF+6JmOsi27/jrysX9MSIryCy8nI1+/QLcF
8i26lAUjxFHfl9lfvua4qZt+uTxF4Vzi0dq/BLEft56wQLRJ0scQy+U+diEkQoPahT4K3qAA84Xq
ci02sKcMTu2eTWAm3GsJyP/ZDFRamnE1DEHvqupV2hJEJj9inM30TKKvvBOk68lgIdg3Bhw8BMzV
zszciMyLUxSoxlOPEvIkQow/xiboWNix6XhqsI+U6oE+hK5wfh36Y1yz1HqodEIGqV7q/fm3tEEw
/LL6VCpsFLzqySvnlLvGfwDBxw3KQLc+mcKgrWlWVNeeGb0iqqqkJ8KIBGvbDvuX5wEv7WSnspfN
3rQ3wD+D9p9rBVVnXe3hH0S2pisH2Al5/2K0j2jwwmnzKG9E027etrH4EmrEsWeAq6z899mHrbO4
bbK0TPYbLWVLJtHL/HKZfZyyWKxLZ74yJWkkaqCmmmEzGyAjUeZCJYj5nCBk5Z+d75WaMEpiaw3k
CAYTQsQY8VpuWNVIY75UwmrcXdiARV+20wz4ZkDJA9TbEj6MqLdS5CezZMuPRV188Y+1ZYTuhhar
FdekNDbMA3bAdgrcW8qxY3jNOMZh7OznKrF65sZRzCVFT20hSRVGrtMDQWf77xe0ieiarou2iEak
XCC6BhT7jZxMB9LMNlF4SeiMO7qVTlcVLQ1v64JqBm6dIojKsJLraXrn8E/EDijslUOGmmht4IcZ
G4Tf7gVjk6jyw+kjvxY4ACNWsSNX6hFqAPjdxNmv9AIY1zKc50FCSFnAb9IhBEvnPqM4L019jB8j
3DZLw2BDvs0NExZJJs23v8NoB2yMkk6FcRiXE3M+4lI54x2ftcn76OgrNYwM6yI9bBx9zSySy1sD
uvpUoWds06An4flhgLeNvsTFyBHsLRqCRuhTWbSKRnZhZFLZs6f4SB9M+g7uc5xYRJDqJvDB3q2X
2Sz3KJnwDeQHqKDH0fPW/cJVEcWsH/6F1rx3ZqRK4n60fU6k5pFJ3XRT4p87ost92mhy95rj7v+z
4Y/O21jdaCceGdVXXPXZyOzpIMXBBOyBettJ0ICRUfJbMsBwHSb/THRYyzQDwwnQvct3ox3TaxHr
sZD8pt1eMitRElpRIGF8Hn4L7zPGdzpEeZ906EbC27xuGtr5Q9fU69ww0fmfMW1DzlM8levF1DiS
aOl4Kv1qFc7MI0g3GtmuYraI21yzqWxVyAmziiF9xP7bTq3dTWi77wId7E9DqktWHEZM28jmD18+
z3QWKn8afhVuiptdckaUeEeXntzw7M2ahs+caGZI+lHOU7IqNJJxSv4GVv/LYSzalgM4Dv8UUUio
alXLS+Nu/5LoTztC70VbQJxEHP9VkHNu+Yg03VZXKltK+C8nU8zL1OfM9flHncbjMjR+1WX8s6DA
iIGP2IyVtt5q2SrLQdlcFWCScnz6IQrVO80IpIMMZNmPosq8h84bwSCEByEZHaeI4oiiyL6ON3rk
aiczGnKZd64fFAjfTgzRP8S8hngOl0GtMoYrwOgal6Zc93CYGmRB31mooK6Xb5b3CDxVs+iFbxrx
vivm1Qw97UZ2z+8JXcspwqgf2occaG9Fk8NMJ79qONWXkimgUoLXl+G2tdGeJFqlpzIWNUbYkIKb
0e4Ku58S0QcEp+j5U6HbjPbhN4Dn72Q23cvDbZRlMruqgNpYWWctKSuBiGvx7mPicg3vDQF5up/i
TiaXHUDO5DAhL6gR2pMud51yDD8NATyAiu9jzoChD4Sp3oPwS0gG2bOGUxRaVTQZKonp6IIBYEm7
KSnfjqp2mdYUEmBpPl2qt19OW5LvWsvqtq1+umbNQ8lsTjPgftH4z6+t0T7rMvwD5Ma/UQVgjYn4
5W2u3OiwfNxefNI0xRxaujMiVXTj/NKwxCxJUwNe1pStrimHtPpYApbUC/DfA4cBA/K4dotT2JGA
aOFnm2WAqpRyH+UZudnqxEhNIKMCjXuGfXz/DgK1AUaAaz8IPD6hYfWBExq8NbSIemPn1bqe7sA2
Yg+XMrZeBt47ORNPhJCvoP8Es5N52O4omvxTiE/Doo3cF5e6Xvs9RimcAdFtWao1QZvWyGzb35If
ySKuz/rlt3vEjuocYGGUFenu+5VxYQhdbYPRz74vfHLi82zj9FVvKy6PTnfwERlJHiIMgJ4se9oi
zu/1RAMCT2RvDbTdFRO09eZV0SCJXmGC/WEoAefD70fEg2KBqv9X4N7akyirbJ+3jVtPRsLlZNy2
8r9kZYNc43y3ykgqww3OvZ1fZJDCBQekjbrJQc0yFQgVYQU2GwejJNXTzAWIZ+vOSlIPlbvCkgV1
dNOCLVY2dhxLT/M+GScxmTmYUG4HZHXseqedUAwQH4tKhy4Y0VoSsmR8EzVrb4wUqNAo/iqMxqyI
24UyHgpVkCNdyICWVEQqiVeCC/s14n7WQL/y9FhMF0eIkh3rN6oRFmI0lc4xxRZHAuJBNuIapw3/
hUYbuYsDIvt7BZDHHG3CsMwwFoJIH/HIALcCpwv3ElNZJoNJ3hoWIoMyEzKa19+nreBsc6CSKAte
uGXKA+CJmAAgYi80sGA9JoOlH1RFCuHJVcPwmg6DJHsLnT3AF8ZPPz2M9I+FRVTU4vDMdTTgFsy/
SHAGdyPw1W1/Bmqdxf9WXfqFwH6NN3H3FZ44JJ12/lRu9YavkPsDBsDuwQ5Jtq7y6XQcyUF7qohE
yhznoQrefFZEv9/Cs6eABnfJrQwYJ9ZwhxwP4a6FZi/Yhh3qh8oLh59ftt6KaXczyGeF3QDLlFLk
OoAhRN38y9fVI/WsB+NMaS0s+KbSWLq9Og7XONmjZCuhL4TGhYvYijmniI72gSD3zVEcRIAj10Mp
2DuLvmj2v8inXSBA+gpYy0bGHJqTzWCgt6q4uqkXXwu/EpS58vmZBKhK46mwjKBlohwCXDEhUUay
YOKYhKsu5kOeUsgQ0VejH3brKne8AR+5U24YtdpybZpyDlPRjIc47Sw7aJA8PmKgfBpYeI05kJBm
PkxGZsY6meP/NCs1ZxWYEUzPqGdI2sXTUvWBLuQVRhsoAM+jb9dYsoa8s3cimBymJJ367gQX04U8
jD7tEWBBORSTGOZxQvI1QnZor1q8+LT1DTkXXutaXBT6OI5KQ7v8IFJkEIlSdVBDfUfHz3MfgUxM
K+/jT9CiT+Fij4aIolABjlx4qN8Yu+oJ2Wg4qBoGfAiM9Kq4S/PmPEYEEdvHlJW66aJ0qdp7gJFS
MB5GJAC2s+6eXI02Ydh/3lnSwXc06BSzfrlOUeImp+OoRPWdmlBJB6RSnH60bT985eq35Xafm5RM
fH54qoxsqphZHbMGOCTepWaAkCef4Cq7EIW+zuo0Y4AtVyI9OBMr2EfF7AWDB51vXLfdUuuMFmvq
7ADLD4XZ++sU7Cz19++vOBFyqnwHqWI7ZSOiquby4hm6CBtSBDkt7EOY7SomleMBDH09NyZ5XDAz
+Sc1FbG9Nqnmp3B1iARkK23jpOQH9uw0B5mNs1ODD20sSdlnbPB8bML6lUSb7I1l2wlTPkl98f/x
xz5aLxPIjkNjlC7ZjmfiRi4ZS9r7Czitk7aiIe/ajqphAb7DAQsYt/+u5jU2XTu/PkpYtic+ghIs
KjrdcH5IRmJJ/XZoeP8tALXG2Jy+C2KOh3Pztl0LxBa8O0WzXyjp6PSU1iO3sXZknWuXqR85W9N0
eW4HDW/jCtwFcPBXk5CgvC0kiQpDuVEroynXe5RSoFm5qE1vTlb/PPsiH3RcSzZ3vukD7qgHepwx
Ko1xEwFnlDwA6pl0wEX9AIlGL/f0BrFtsCquWFQUf9zNKrk0O4sk+Tqc8Lfh98Lc9TjXef8eJ5aZ
wtIX4hZKyg5/JgMF9P0LDwymm9+tO+6u+oSagpuWJEXHpi+pel01LvY6IfbAThDQTbyq9kLoLLNg
R0bQiONjRqu4WjsnpSZdwNwLZnq1sWn3PcfD8o/B8KpQrUVRiML2KUccK8p/1dg5tAHDJ4z80Dfd
boKDvBYlraqQci9djQDZrbIpXb+829Bu/bHJ04f/Vv7lAPki/0PRisyHesM0C0RAn+mZRN6oHDPa
9QY0dFJ954rJLxDmwluvX/HZDJTewUpbOSVyTKnJ14cu4QN/cdiBeDqHOu385xxjmyfreFtJFmsN
IoacX2rso0ScY6QfjAXKOm/7GzxQnVz+AnJcmPQH/IBLOrV1b3U9WYWfBFXoLVRXSwlySthdeFix
JjYZFgU9cWDPy8MHyZ8FjGD+PV903WNASf7tx4hapzvxeOvxT18J3lrd1RUY2ik4kzk/CVaIVVSa
3VpXWy+BPialyFg9judSu6IB5Ywys9YXzvaPomLiCWKCYHpwFsifSSlNR4tA+ejEpMGjeZBuYvNm
PBlFMZY3QRn3g5y40PBJpRp+aRq4I4YY+LEIpcb4j19hXj0h8TplCyycnd4K7i9pXwnPO9tumcJQ
4QZMkWalchkA2rxiWAVLk+33YRbQI8FXyVfpFbdo+bjk4SxhKztdaaUQpiUDsb57H+x2rA0YCyiN
3F4kvxksuRZAw5vtsLTAEhDaitaYLWLJbJspgzIl5X9b6NP/Ok0YlN4A/+nY/A+HfV5xqFW1j3Xa
02k7KuDWzRqJQauPyQKcly1xgFlawZe92Xjm4k9EX5sp8pONpqerm7rtfMM8qlcSJ8kmhMesHXw7
9uE6vJywoP/2viyRRX1wVaks2WC/bFmMrvc+XicQCqbU0jG/qDgguUoYLjYypaXpj+mCjqd9xSuw
3RUiEfnHohQYylrl83Lw6vdZI3z0v2eOJC612avWVzRkjqV+1556KgZnj5aUaFJy9HdFNCk26wJu
o7iRrgwG/nskHmZdRIKmINT/MQr0eX6BgTS4zTpSG6gA0d6tPuZMDko+eKageVE0pfMyNWyRMwBG
OtHgN3GphLkr+Futotqq1GfPwOnENclfbeoaardr7HMFzjYkhUbiCX5LU2SQj97pqXfdTGu/r8Vb
dwXjxcofAB68Eaotz3AdTHG04nBwp79Gkpx6QHIV2zlOTYMohnTgstpRYTK2sKBC4IEKVspPMD/Q
+xDhtx7rzk9Nm/zw867H5lRq+Z5TK73GSl/ekI4l7uASrpCIPgqgIqf3dBL8phVIbPwEff59mQnM
DTRJvKboqrFIRQ9nNSbOFs/+8Q/VGvz7UTHrIO2PJvToL1cRcxwZda7tbwHCLLwdiyM7UjWi191S
pkRePC0BwZC1d98QiRPbNTYBB9odKamkE9JN6XMlvywAiV0zz55lvoSzK3NSqIGI7mOL0q2oBDqO
SsIYBm3at2vYD55YB5BK9rIozr33NF1sXtFRdLtwL1p0cf9MVvCsKJ8ArPjabd8K0PnYZ/N6YytO
LSb3whna5xMYy3AA/m51hqXMoOQEdms8PLWLqeyTX1cWYB/03qoaDXADp4z7pNX5xiRG+KVKzXCP
F+VqRPPXkq3A0todE+1Xo0PCwm94jVVUFz6qRXNNOb19h15Qg3bT+GMl4ycAU7sQCKbdSjofr4s/
30aOvWM77FzZwgX3VFGfCOHGVIMRLy+ycoHndEza+RrrCVI24tIwTsFx+tNS/A+M78Fl0KTBBcJr
9SgZC8bVxSHrWapmL46nYvGsugzCLPI5Q0hQHRCo0kuH9ntl9mBDSzs+ozPRDuSeTsLjZIkkGpDD
lzmkTPbDHoufgwyOjzb1iDH35QsMgVRifMR7xL+NBS4OhCugneBGVNFrqp0u9a4M2OFZlBFkq7+B
4UfwvQGpPOotZzawNeFPrHCwOeQ+CAJn6IhTB/EljLLlXVIjdflkOITQW6kg9nKmbK2rLl6dyLqD
UxSZLgGsXTMU7LS4KU5nZzdcFT+OZSSYqFPvGZ9oR6lBMOq+xaO7W6tmvZaLcJhYi5pzfq6wZeo4
aJVP1GdA4Rbk6lRCovorOKJtuOL4HqG4raACgX8n/f14a2XcOK8JmkdcBkgjA4zrq/nlH4EKi2PE
r64jfPwlrfX//I/cFe2l1IsaoxFqxokYVICqJn+ht9UnYA4X6hdFMFpnJ2X8Jv7bXcSxFu1n07n6
X6UZXmUbUUaQaxEd8ArJK+3fSCvxwbVRlbakWbtTdRVt4RTuPyGm/trLF+MDE/0ihm2C15n6m+BR
4TNd8QIPNArCtI2EKZIR7HCMY3i1g28zcMRA0qtCYtZGTDmtUzN2iZ6GVI/Gof9QIcHePvMqydzi
RTMVtCXnzQEYKLQTSq1NgOKeRbD2/T6/gf+Kd1Zdafp1Z4H5LDObUR6I1D9fUawGAmSG3CXLQveo
PVHo4NZzkxwWJ/7CHf86Kp5I4Pwes78CQfqjjQjxXGI1j7vTscyjOBKcg60E3Yw4ehoNA7KXMSqp
x3CiRfz96uORC0YHYr/RpvM1ofOa1L7UtK6Np2Wdn5vScVnktPYiltAnAekeGauCNzEHTwYeqHXr
9hM8Bm1QU3UyJy4Mdd+nJ49+ObXgndr5TYWrpblD3GHI1XSpNMS7MW+SslEGPnlYDAvFFRbYDTlZ
5gCrEbgGDtW6k4ydrYkG/o+UspIKowUPzCmlsASDxgCOusUhWYAdH7RXZs73gGn1d74IFdtwkygK
nkWldHSuZqL191Z+ywajlrsgSG0rKnmJR5zhslwYFeLPL2eb9ofT4CLbe66sNAeSnBQQufisgC4m
1s2ug0iH2gRVN9Vve3IAHOxuoHJiVzFc2KJaPEuGPupho3xI/7XtOE+2ze1CsMhKdbsm1VqQwTvb
JqiTbnzqhypae7+qhTUjCdj5BxxdCmi1cIWR2eKDDayvm8//DBG3Mv3/TUVnNhTRvGoUS+gYIgVm
BiVByuQpDpO7U6mKYkEk1o0+RxxhnsSm5v3psGbnP2CDQ0ALUYKMMlK/ZiLxw4OkWvLxZw+G8vEg
yQqBA7yj8paH9kHMXjjRfWSOgJRn0cwayqSJ9fqkYOVTPELCC6kgx6z4DPUoPe4kJfnQ6gieS1tG
27Cg513BSAziw0Md2nLxq7dKJWMzd8HsuEAUCHrYw1GrkXaq4eu7a/ulRxhRel/+3NHgKJpze4oE
Hu7nolvE8NZSZB7eJci08lEPLytpMIvvA2utvHS7HpYamrnbs72Hb3uyohkuKhh2domNXfTU4v7J
WOFp94yTmOY4gYXz32mbzOuG9WX0pFa27Zj2VRsgLKfUVF8AvSJdWrLViVrSU8AiEl8crBJyQDwn
1vWWe40VUfaRT4VKc3/mY+LTqDsaYqWvmGdCKfyVwFfI+dQV/kMf3hDfoNvJqvUdwHSwX17KhZt5
i4droUV+XNPuYZ5q+As2DeniZZS1viHxGvKcCM84Dh/uRrzYgPxkfdF5Z9wED9IefPj/asSlms5s
jH4RQ2CL/H/YLe/rndyAk/d4KHTTOw5i5BfvgcKKz/01i8L2fLpM5BpXzXIX3C5cuypeJF6aeOQj
AMcQ5eqY7f5hnXx8r7NSV71QJH75qpuw0X2iKMTQ/vgYhrSU8jwPyAVafPQAanzfcmvozxOFcqST
qhG++QHWS7sXgaSbBqTmcq02dWiHt0Ect2M0Opx6jRpanEPHEOmvI8XIomjZ7xxG2U/MzNBjJJTO
+G9Rq6OkTiEd27cIAHU9zgHEukhyymO3JZdn4Nt2q3/DcrrBLZ9jmsT+fLUzBCHL4WLrTmzP1ATC
2obafLRlTYIiICKDxq0YtfDWDHBMFwsP573HdpLOhHIJMqULqUEU3sgsUFQXSPNAmTLzX6/fMPON
9EcVCqIMg6kbda/bILVBdHUm5Q/4WBnttZJtFOrTm67K/nsU1EpeqFkOcwqQp77jYDDwSdyLXxt+
Z7EGkXbGsL30Z5woGVCYX3RlDlHTISk9IzwQEm9RV2P2nPmUctJ+fQL+EH76cMQ0bAmBmrUVebEg
TKh//Uu1nNhU0gFnEo+EHDZjpDJFyuXepNoet0gam1QYQ88YVQtxi7BdbBDjZBe7RAQYQMkuS1Ry
K0cK2gMzIG5/vQzCcyCrjwZw9LFeX6Gh0wsNO82uMkFJSBco5Z4bGk7W+3pmwgWEwMkKtlqDCycV
yBk7rgoYm2HPutto/w5tDHmdLv4D/+a5quxojKHURuFyrqQQKUtUxIJy7FwmY6y5iJAJtdKKtFKh
yFtNO0fS951yakpSc8Ixm/LtGlCYm6vUXZC5c2r07CGHBpV+k6wpO4b9j3CGfVKxPyWi3CaSjxLb
ppk9JajAtS9YQC1OjX9oRCUQVvWtbxwaELkCmCX8lt0uN29DH6TKzj+Vk8hDjvObI+Egi95nH8hE
HTmVEGdPBtTZcrfR+MJ9Wo4mP9PlVHUHDi6is/8mo2e+JUWfoAgnuLegUzZM4/j+yndl1FBFZyzW
Pw3kjbH1c/3e/YRW0kCiP9mY5vNJCWmgPksOox3ENYPlO0cSI2swDvWU4ooe5Pme/Y5QJaqxQ75z
TqGIvoIl8+euMPppIl31wiylPV+n9v65eKwccsZSX6N+98yoQErbUNk42R7v5AJVH4ZuM3XW4KPe
HuLwh5F0WB9Mth95mzxEbU0XgRNzg5eGfS27JSCIjHyNRjesHGTlHOHXCSm1tjHpqfKjk8okA56T
se7/prgackfXg5wZK4ObcxhGM47XP6VZZnb3dXBA85pffvoOdv2tJA3JTj6uY+050y93yaVBp15v
sv5VHFHr121/H9pMtuXM9hgajySVB3FicXxL1+T2LkNZfW89y5BXG4G1EzcCJhuBJvXzJn09MZzE
Jy/+tYNsNjl/QP7j3Cjec1SagsdMl7NREkFaiBW6EijxKPznyJy546Zo5ZqfczLTacKTbFgrPZwW
7Ebm/H6GWq1pWvQGVlRHlf/HYH/EiEPy8Av8lcoptUQMoMG3UjeV+lt6wVFZLWKEKCuNpoAM9HhK
hSlGXcguf6tMvxyCoDKG+c6aV7ubBhTc6jbNLjPhgvWSdc/Y0k0rGo1/kE4pTol/NdX48d95AYOn
Xqa+XcMqRgjYla7E0pUqymT+uZCwEXd6N6nNTKyJg7uGda1DVikecjLMifSi2xXWd1EzQRDPcT84
bjW2N1wPMQZAf6Cf40Ryz4kv3Uh+491zid7uFK/cBk2B1XKUQ2SsC3tcGVz9q3rRhzckqWK3TMVN
1QrNFTVEDcolUrxkH9CAhxeQQAcGpzVyDy4FYJ5Wrn8vxjDAMPTXmGE/EycffoytaRVr2S6yojio
N6R9V7xHO50Eek3+nQAdcC1utao/QM4A7z4wx8iaaieTfF4qHEcJYzJSz/vSHYfPyh1jIFpo9wRD
dTTUvi/kD2P+x+X9YF4fwDHnMm22o9vs3snQCApoUi5/QjYnQQhusCCF2D55zlTS12ZaPG0G1F3G
KTovF280jrbslqZ5wYUDJA5xxIl0nzTwSSPIqUEd8gDRL1Atist9KqhFfBLSn6LrGkQU7nFTUFDP
lfmXSiJRLii2fJzf5+ndApDwrnQfG7XUMNaKo5QIXPEtDv56hlO3CXm090llqAIJJxopn06BI7uV
YxFAaaEzyB/naxURbyCG3I1FAm7FahnZADCvMJ78lcurgg6fvBKhiq9GogMzz+uMwa2Emfsa1+lm
X85EW9CwVHjvAFYwIoe39bBGy5KYleLgw01bcEHJlSEVwE7WBn+v+QtXaszZQ4qIQ3MutYzKhzg/
rFU92qZDbtJsHhztpjkAO8srEjIB3eYaASOM1VzQlh7WaQNXd+7RkCuTQ9282lrKKGr6YmscBo3i
mxu5jYC1/xbiZudl5EhPJrTzaTNCZgk4F+Qjvxfsl0DrPE0qJrqtMdooWfkOKZwqDfPOIb1R27+i
zeJqaPkXjx/2IGAJ+VQJszLV0ryS8p9aofgAyyr8iz/mneRoLyL/+CMPCOT4CCnZux4yEqH2lrgU
TI4M5eOPVAffzUqMnHSnHyB0OH6jiC6SnGAb1WxhD6obfYb3lJ5+7R7W8iHnbW/+EDwZSI61zJcI
XlcIe6MaC1YAzlcD367bzjHnzfnAfqdKlBmMcP9reMjJWipzHbjh+HgBv6E9szUf2YFf+OeGuhaT
AcZgnZ3NbxDX6VAdJlE8DgA+LrRKhACW9Qz2yLXYikWeP9SkfFSki9uvhv/kUBJ/lF8nz9cjaUHo
hCk2MVl7jTt3f6Itd4UvZNaJDNolq91kOOsgQG2eegfn5F73lmC/eUdnvH4TFXCyeIm+igI0nHDw
LjTP9t7/VREQEv/FZgbdvUvn5510JQdg/Pa5xDaAatCf70xe8XFauiMPW/00KbdMkhdmFBlubiYf
ZcPt9KM5m6wW9783HqF4nhvKYDyZyduFVnXdhl/EV1b40YElVc/TRdneMiQkYb1zOGpgM/h636Gt
WaEArYKA2wVXhIR9mHhtKfkks+zBD6q6znpt1QgCQbiqURQY7rDegk8MKRRWnLEUkOlp1c8wB/wI
4GS3uLmJl+PytrTIw04UKF58EtjL5WznN0OkuRbsHZ8KlqYU8phgSofi6CFNyYHuO9ZXII9+ADZB
czh37n3+8sY9pCYeW3t5LjH0LW/uQnKELNQ4mfN0zFmRqLX8NQ5fmcllOT42wIrwwbCqCJ7xAa/u
SHSCrnhaYWN9AhgSdgp/szEsPqLKxD8nzVp6+rhYWIqxpKRnRmKmw3Un1AvbBh8KUI+xR9K08bzL
LKBIVZ3FbrbG8aeR7QZdNLLYs9jEKqlaWWjiLejDO2tO/bwypvou3OmLPXQqMFA8gG2Tr4gY0YPS
CjNhQTxNonQBeZmUVy47u4Os6jbalybq1s9Rl6pER25b0NrsDGhDlGPP36FNWBQphLxLAo/sozoG
8PDNrT/ywWyRvf4zFqv10CmgOknp1dbrlodAEerwrLvCE7w/ZOfvP5mxPWv30+eAbHuCnySw+ey6
MYZoDYWPlKqS2YYwFHNMoBXTSjXpR/+TZ79EHvO1RYrSl5bEb4Uwypey2xw8ZnqCKdWJUrkf131H
wNGmZ5qpiTsgHScNi3jSEvu0+zukEk6gAkM3gRlGJqMFH4+DffzcYW5jTfpMVtyKmukw2GKUhQi0
nX4/ySwTsN0UkzjUzb7X+oMqYQutELlILmoFGVUjru5/O1adjLFgRAceymui46p/mNRy6mlKN64T
HSRRYxVjUoqsBq+rLWR3hjc92cpSmdUdYh3a+URercJ6QKZVKcLWjnegvm9JD4lhD09VJXcvAq+z
eHigfE6bPMYEU2U/sPL7mXk5Gf0Z02mPe8IentcNF/oKyUBoEuBPOaALgwrsR/R+CSYZMtLfjcl4
dDXskb3G3u1SxVCXZ6wEHCZY2z3RV8FDI1CURYL40Zn2DvLFdvHD698xteZxPMWVK1PVNLloh26D
afKZJKcRzi+Sr0vYzrha4payWv5/I/S6+ilnFqrcWDgrmwFPxoyXZj31cNsEOwH5DBE7Ky1lSIEX
irKqNIWZ8/jGFPCSNqNwu2gKue1KZgkB8g/5LCJxHrZ4rNw2dir7wq0hSaRmoyQ7ZwpyBtrGxnos
KdcUrzz6yTX5h5GUAW+wiUc6uEtLXWxXl/jOy3mY/sqRL37H9hv8S3xQ3CsAviHoDd9N3OPOdwRT
T0b6VT//PpNLBKU6QORGqs7RnP5BFJ53DeQvis1YS+rmvphecWjyAtGcINMJ9SwtdXEln2EjT0SD
AgpoblhOA5AuNv2qeuwU11ape5/N8pOqBDGc9cYeOVioAWdZYhuRipV5ti2habkNC1jIBmsNvnjj
CxOWmj0HA7phUt1YP5gxEm3Fnj0C0HNCnD+bx9grRKX0ECXt7JIoOy1rg+LwxwwBwDD9Ai7p3+1+
ZVqauo2iYyKzaV9XkRrGKxu0qs+oermlJa4XlwwRv0hg3rfS2xIG37+384vQYOX0cabitbohpXB+
M/dYP8qAdr8qWblGwioi38369EdU86L9YENXi8HW+du8U4XxuBI3+Wm9+j23/jpEi76Zr6U9go63
XEURP7+JrorKOqUFbeGsy279JkVCxYFUt6M/SBUn72WtYZnC0+50I6Ugd4pDqbNjKBulJhQshe0V
dyRa1jwO82paC8MOZcMhnbGGbppWN3pp4SfO+gsaWAWNNhMMwZqriCIcNQ2l6V7WfvVFvwEWA/yx
xjPPpcBm+b7gVCd7/Mahw2iKZuBUPh9u3LRTzLywwXZ1FoNgwwMDyweUpNQTIAVssaJi8PnFPARM
pDSoqF+/oiJJjswxqDHD2ES7ROCIHZTqk4wEB5/RJQk8nUtOwIdxKnKukysvFRR3W1j9sAEy6wwz
ZRrKNxd43eV3IU2JMbjK8k6EdNYti+sDbS93BWls64sbxlWnw8nge5gCbBVQA00slaqFk5IQRNkW
LUlPtA5kcL8uj5Lf/x2WNy/fuLGsgmmfX1MuH8jGu8+b83JRAeTUhbTrJrE3lPeLKNGuypaYg0t1
LlL86jvV63cVZJASCZutYF3q6AS1VuXcf3uVqanerHBerDA72nw3acJ4pk7T1dXUF+CigW2zcg0E
vTjo/CqL2mGlq1/L5JfmRzo9TkEgFWHGoLkgRwnOB9ecF5DTJp0XK1kE+/2hsdRBrDoytDUwPgh7
/QGRvkORpeYaix1QuYTFpWcM709Mw7BLJLqFuyMMXJLqF+OM1FEZt4E2BtnT/WHvfi5kmJWpkawi
iYnUvwFj7N3udCMGIm4HoUcazix6EHOB8SqF/5GBd0EpyJpuvwakl+Zp0CRUPZRtNnmNZPjhdGTd
Tt6ZehyMNxxGVZEmMIulXbXRkgen7sRgdMVRmQqgElIEepuL+kxsFJBwoi3RHLssmLiF6vPqpTHx
QBRtOBVvtUAPm+VDy38tC/jrqZpim+ideeKkIrM1ZgY1rSWBHru8z5D0Bf91MgJuvh1T4EDbGLIx
/FZMlincpCFlvrpkGFSbhe+x6E/1iiUmhc1XLYiB7jTFkmMuX9/vqRENJkxr6KCpybyWazuHv2rM
3pjuZ3JPJrRHv+tvpx0UgKEblCkAATEOatK4Si4rfexa/S0KrRpFz17ClNbxPDVsEykZzB6ntKeO
xLeA/fTRZHqJTOqq3h6rgDnz831sCe0hRNQ/tqqLBRKrZS6bgzZO6w5B8S9cmHf2U1jX4fttIG4+
3NLp3ggNnhu31wPkl9HSUm70NMDwSTfTXQHbv8359bLIViFw6z4Zgbsha9i34tyww/cmawxVxmz/
e5/JtWzwPXuHVy79rpHRIV02qdyeC+FCrvQCeA5dpHUKwuS1LqLRxeN4hwrGAQAz8lfwXIgw4XMq
AyXyluEECqEZcz+s76ySvIs2reiGo0ZHuwPVH4h6DhSZQDmwYJ8rHn3Su27yZAFCFIdgT/g7zUzs
9kjIaZleo5HzgVhM9CWSfBnt1XYNJKaM+pFI/J1K9He1c5Gyv6i16OmPtGsWegp+pxQqrSrkLiw3
aSMpcifmTsnXKp3JvKPgQtlwb3bLkWSYtxmxI72EBMALQGasmUSzqgjEqxXUXkItj5pbEmYCuINW
SaAWZclqTn/TI49mTT4l4tMQGfUATsLJ5vjwGmHpvsxU7eSVkHlQZMST4/V6i7vOBanMoq3UelQE
6aGxzToPdZ157nd4B93pLMw0VINgzxeuh5zv1hPxxy2DXcblwd4zR0DEkjoBweFWyu2+P7kF3GjN
7kVz11JiBSPm/Ehpu2+Vor5iP+lzTwOiSSWsRf3JvP/UTqACkyGkAK8cHDJo1JvLqSOYXlthHjKj
Ixdny65QnVl2DvYfe3UhsJsb3FcU68nnqpi8JHHX+XBMaLQwC+fmWB+iO/ZHc8h7QafrqA5x4y2m
3FYa3l6NZzl65hU4ihDyNRAsyAooTRmcNjFmsM3FiHd7VJkwmSozqQ0/Y3H9ncOMU44fBBAlH8UV
nharlzLfhDXBAm8s7dax+L5Ejtw/fBoBhfU5N94ykUwoWMlzIh80jrPSf39UZ5Nc0LWKFLGLFhXe
qIkqo6IdIpR7Ls1b1j1M6oOW4fNn3ZgUtUrn8mvbzqte7AkmpKbgP3E/qrPunngYhpotweEVlK6o
GsrnbvvyN/8CtknPmL4sUv2AM3qUYg0xrODDuQqWN4B++TNiez3oO7yovj6V7Ya2XRBh4siEnn7r
vQNpC8IJLWEC2xrk36PZvb41lDECHi7OLHaWLmyG8/RlHvoOW/7KVp2J6j4nFRJ/x7PVPWOlvfvd
7Q4yMf/k6TU+O2cBuCQvlhFqR1dGel+F56RQHDtxHX8HZBHdr+YGfHeymo5zaSdXU2hmTGqW5JVb
6SXxUbozzPG6kNUd0nb7fxRnI3zoOX/6yQT0aVv6/TIH/5xnIYcT9oeNPGdLm5YgnvSAQt/BtQdI
m3haSqV3qkr9A5fH2DOIonRV6ujHCuYlPrEQc3ceDj60Hl6ZIOJB+/aQXQH8NH8Q12nxKw6xktCp
ex0YzdRpV/KGMTm984CeeyuqQcEeajHVbssbPQzdNFrhHmTQ99ykpZhB7LMG8u6ekSTHPIhl64XJ
sAMYd2oDWY+qVU9XYRpnBK9unobxt32kHq9f6X6r4g8c4+kYUpxWuXPM8uhYtm7FlnxBUu266m90
mIDApxpup4CaNErQJfFCMwSXN2ELej7KkyLI+NyO557+L+cwMgdiK8yg2RW/zPF2v52Wx+YcD2lV
iCMQzRa67rqPpSSNwud0NfMwsAeIen85+FPGvYsqwFvcsSFVlRnTSyQi4CbV2o1S6Et2O/cPzqxB
vYbMS116ZJzQDquoh6oQtHKEaZEGPHRUjouUE+ik+ArbJRJ53DiPg85W7XfaySYDCUoXonTnsBa8
QrVLzq2FLJ9p2EyUysobUCafGC4W23vcrSrvE7XsQX4vEbhr7YfDBA91Ua2fzzKtr9UYG7OTI83h
yBaaVQ7rJGCefmPQUPFsxE0XMNWn0j4tIzGbvO8WoS7SVhHzgd+JmI5xobUooP0tJq9fHfb4PLBf
OuFxGgcR+48Ahx2+/n8dqsZksyGmJNk5t27dXWg3duhn98DjmVUmyBCOWV1qQcVGLwoUXJKBpuFt
s0ovafsFj2JZkZYUmHQLv6ydgxJoO5o/umx4tV3UINevCAKM+4gb31vx33LzyumqTQBcBV2Da8qx
u8K7oMRRsDz+UkFZBkEZ7mwlbvAQksPbpsj2izFa2Ce3UBJxbJIB22rGepbKNWJ8heF/tDfVtNjK
npd8lDkRLq0Ss3lWyfRV7ZDKOOprajSzRmGdpAgPu0JNMb8gTzXpoAunaX4G7OgfDhBvnjnjVgJA
iPVvhE3dOTmyIGGUglEniaPO8mRglPSz7pHkoDMpspP41kGisSs9q0wUZYa3eK6llV6ptfXRgq9m
vcupPsjUkEBmqJadpj/DvFWg5+kdKKrBoVvwPxO//oOpLARAPYI12MQKRJpkAo9tiEyB4kU9VXqG
j3bX91KCK5WXWrviCXRt0XWi5YE7XfA+wKkIhE58fqWVdj+WyaS2P++cf3Myx7iwsgn8LAbGBDqH
Exi2MeTmR0T204F8Xo8IJhajqpkGhYBqzZcELXN8jO36fb3ywYbvd7S4pJu1PPeukzYgd3GVzkmu
ObI8Viub93sCA0A2HeE6GfS4NoEE/OkcGe0dhsIuzZRQ7UXeXAqrvxNUd2JYuuFZno9AmWVrZsUb
xP7ZszScGiqA4U4y4DeL57sv/V6Ltaeun1fF2gsvO9CazsoRqlOCOHLhTGeyqo9b6XdpfI9K8g4B
7fK3aSzfL2jIXtbMgWueogKcmiAWhVoRY4ycFK7AB7T6TjAWP5MOKhIPLOKH151xyTaVkrYhXWQg
sLKwUhDmLnDCIUN5J09FEgyZki6wHRCqMT4q1dI20duNIQbPpqL4SJKjUbBgAHEY/tS9fiTIhQrC
4hDtadyjGjl8JzFWf77xnp4jkNXd/ofAlKhaamR0NXOHKZIh6uxGmXjEwo8Ev0ixIqaYbh2hc5y5
IqUL++HP/f6Mfexo35BB4p2/fPYtSBOIgHrzVBpdzSO05mYndPIgkddJaFlv+YoUez7nc1xziXJC
apVKzau1IWoDhGAUIkDB/WzYPnPViVOSizon90RObJj5OuQrfqBAKCYHfxqnvhYJIbZSU7DvVifp
NdA2UF7StRlhsEVDl2W5zUIci2rVT/TOGDh6kQeHsHZX7/gkI9qoqbAFlAoUDycoFjDsoq4aKxT0
YWMG7Jbmqdjl3gpB1vTLkGU0i/f4VQyYnI9NSfCd5/FQBGBO6EPsmCLvonXTA3yoba3HAWQK/JyK
lqHoxx0GAp8VqDM2IJFM6v+c3T5BZZSWaLQ3wGmMB7sK9WElf568Tesg/oFobvFJrq35tHf4pR9I
xOTGLEhFFPQRjyAZkPQD7tlnYWUK8a//4qIpoSgqkoKbWEznJcdXcEdhFxA1/Imlm3UNgIsBeUlM
zwBASXrb7rCu+JN4oOpzwQnAhTOH7kOrzY9DpvHEokOUivlZocmdfcwmtp2otFOA8cLDG9MM4LUZ
PVismRKlc/gbSuqldhp4EjWM2DL6LTDagFtw0Tftl5np/tsQvML5+GAKtQythrWTJyft3dbivJXw
0haTIfEOfVDjlntg29SJSk9ja8UMNrb9jqP6t3t3VVynX758ECmG3f2vl5GJ2pUusxhe1owQMlc7
WRdAEQQP9/DBLLm+e3YwwMLZ1YerwXN3zn4mFs5CQnglGvoUVwrskNlJg6TInVVl4R44wpchNBum
9ddta0AOyFk+w4TT3RzSWkoKgX+UwAOVnW44hDn/44/XyU+GdTN4U4tWEOk0uOByEMzUl0RUxrDo
8NG6gdWZuSYy1pXSMEPVR7+ZzeuT0HiZlr5pBUyX3gFTsI70T9tOv5c3mSSltnci1AAJsDNsUI+i
i3BpNGs50o42bcgttYKk/Tz7nuSTdytdnAJ4jBGIR5SkLqHMXAfttTgGq1NxH+ZUqdaYXBeb4oDw
yJvjnSZKJ8Nb4rMIQUutJBvLkseDxjGBiJiXgIbc7OmpdGR9vTAmbHGgxhhz3YUO0nGrh4D6BpQs
bUH8CMNRbxomA2WyFUFB2cBSdAOo0MrHsSHVJhhnbW/+k2QAM38GvKF4zA6iZ4eX9J9auJufWxvf
q1iwN0QTQ4POvsLnhB5FL/2ugMCnVQ6gZLckPtBDSFwEo2FuLzGT6KYDTPEdWyVZrcNglDHjeoCM
ag1ufdO5Cx0elXktXTLK3cLrzT6XHZoHNjlMLZkZoA2BimweE4/a8N45+/yng81dL1bCp5pZfy9M
xWdhr/VxBWiKJ8WsDLb8K9aFbnlBNMqZrtuyOhXhuBrvm06sYwEYq643Pi5KxXnTLjYWCPNVH01l
la/VxPkrdmwnZN9h1XZjHC6JWfXeSQ/7hR49fVu6IzSxJtPljhXiwjEEU2StrPs1wRd/3brN3gyU
WqxS7IdA5HWcK3JqPEARRllXNYCGs1zb1Rit9HxiN3Q3kxqLnKZtkGERR++uACpncqeqbSzvcrP2
gOhnKwnP3OF6QEdAtjNQX6kCTO+isO2+U3MWnTT62fG88tBkryS7zI+KfuwGE4vM731xU+LofcWh
aLo3GXUeuYU6E+2addgGVq2CRausaaT0LWSYDJbpdDOXJxGvrczSU6Jk6+Vm+B/X/WaVCEon+/UM
T1u6/0lng1G2XWPM9+ERVcortN1E37d/Rk/ZXnsMb4/Z9tEpRcy40dM5Qhs54LjcYqmq9kCvoY1e
ujDp4RPBqYPkiB9Jln+PNJsmeB3CpBKRMrLonmI393df6aupaMQsj3yh39RdpCYqOwsRwbfYytgZ
eDxC6zU8MI5TwINTdfgCgS1gX8KdD4YNMMRZHevm8F/ZMR2afh2W+5BIZ7khUF8nHxuHUqAF/e33
V/Ysq+svgkARvbdTtYAZLawpZi9Ytcd1A3PDX0erLVuK6K8TF4GymmmF/ksCsHtQN7C0BC2r2Hej
0oXRBejXQZh8GK9WbWnejrrI/Nw7cOH3RnJuGIV1k16oWbKXdrCLvO7J6Ahf8ZKM3CstTAd5NupG
uhEqjl2KMWZV2gLvY3iXIqHB4R12hErEFADHnhp0rw1PbrSOI07LKJcanSJy9lvpd/oiTNr7V3/B
DWfSR3CQ8dnb7SM/fIhfalE/khClndd5FEhEzr/MBtbXpYvg4c7PVWS6lwoo7mTFrx4AwfLYR7GL
AxDuisksDNw3GEiF6f6tpBo1OYKQVKcK/C+B+IqSNlBO3dXJNhok9+HcpIbrNvTJm7NA5kI8/ozi
o1+6qgSFbhDCxP3CM2Y3tlA6uS3Rc0s/j0vgJIOs2gT1qNJjZ2+pCz4USuK+UtJ763pp2Rjlw52I
43b+soTXHdcdvO464JlWrEc55kaObio6Vs4qnySa3MAqY3EQSpST3ofUMXXheDITPtLfCKEH/W0S
S/GZNQcrFFKAUhoZKEyIwO8aJobJ1WEANVL1RYPkAzK7IgoFnAHjJfGeqacYsErbQOTSvgq+XM/Z
8tO7T8jMDw7TQYlQJDUXvhpY/L/6pT4DwWvbzqQZj+/KLajtOB1M1L9MDLcLenoCMIDL1w1S9bkL
IR16ajFE9+B9QFexWSZP1sGRhWoDRCxEi9nPpmwQdbImdFivG2b40of45SxJP6l++5J0OJn0RIkA
px4FEK6i12MSAylQUHN4+VJ+nb58sClQvT5laj17TI4LzrwQmDbLawdv2s4ugJ2giXOAkDiqMcPL
xVV2dIBhkgiQv/Rrd5qtWU/YWcIaqnFqfKX5M2jQ2kQnwfgIbff68m3mgpDJq9bZWk29krmrqXf2
OLPIadRv5cfL8nN/pTJ/OaLQlw47SrOk0kq3yWtiYYNK7HxuuZd2nNnoLISYz7RYpXrflqmL/QNM
bVOdWNQJlr20lDY5vmDYyG14yW6xuJgD9xOhF4YbPVtdQPkhfytL/umpaNvwqplrY2qDjat4wqFx
XtSVqgBTOb0NYPzcuriHnnvzQDa1FGiGm9W5KvjU8giuJ1oo9zb/C3ffBeMr7IY8twLnRFuTH8KT
/JOkMdotLnXiMuja5UJv80W6ADt3QhKChiT9gZYpd6jorebsdlwdjhrZjUjAtzEh9XQIV/DWKXLJ
wZIy+gd/gv5emkMt2tqdNBbXTsYLeKRIROh9KirJBFfRQ0ckhUqDUAF2UwgjXIyxGW3LumEqNBzb
DZ3Bfs6K5emSTRqjz7pAqhNY6FbqhOGUJtde6RgCtAUxmRNf4MJb9/7hReFb57TIKBkl8zyufUsy
1DOxQjoSwoWjzWccMJ0ULu0rhI9XFbzkGv/WSkud3fvkajILxi3+rBdVygb4TZKc8o/AKpTYiZHM
q43Nc2liPKEcUZQlNv9NwIZJySEEbt9CVu9XMS7hoChHaS+NbJYm52mqRAFWSh0VZVdHWiB8ToQ+
9EuDMOAjR3KuMgsjIlEAr5zpOI09fSRfQt4B7c4rvbrIUoAh+iCH7ugrUr6PL0etaOI2BgrE1ejm
r4Eb2eAyYZ8m/cLQqa7/1WBaxxA9HWyhZvbEdMtjeusW8BZFP4JC0E/BMn3cd5kjlN/fbLqIxyWF
8anwRNAHx3XB/tA3iUzrfC/CllyI9hufzexTFDi9oNOBVgzHYg5ASlkvZco9SWEvhVrHgEamGYs6
NxNJ5Tte9O2IrDEzGGjE1s/LN6xXHA+qs7/aRhtoGvHQju5ON0jNKOy68FSZgqBrG+85pm9bzXDu
1B/v+j1UO2ag2DokOj0fxKpFYIq6TQ/UPhzWPGOhA2dV1vw6fY0w7tJSB/cA9WxypMWsuEfqAwRA
zTCIGcU8Yi5zGyzQ2n+NE9iGNk/KVrHrozidsvrSffYp/n78gGYXzJExdDscBqq0wXOvS5skHStk
x5Bw/EcQwCeTV3iWTNIAh85bjoO9S4LgR80UX7faIt/95C27nZ/4C+sz8SaJR/i1vRF2gWcPXNmw
F1H7+gxemzZixv9eBZ2S7SA6OUbdfaTyTH0bhei+qeQy9Ik5zGm2tH7/QzPVtMDH/q8aZm4Kl/IV
zIxPy+UEDU6C/5uySNdBjZSER4GTjgagFDLkfreUIPEEy1UEjFwg4mrp9YAASZpyHicw5f+Ext0x
SkbGnllwietXXx4fa7RMl79Ny0W/s0yuCHiEF/3e5FazzdZe5aTEydKOdRQf7MYrWjXz9iFTi9HS
0x2Lo7yr5QfcqiYdB9LIG9HBNLuqsV9Z8WM3jxUM2Za255db1sVHzM3hWvcIflPx3fCcpZZ1TBRm
Tiw21eUmudsPBTCx8kJSanPdEFxynV4Pg9NswBOzOeRmx0o9wfRvspF1PZrIF6dfA1MA3gEVS3pS
MwSElbMz8nU2y+f6aK/otg6FuqtyJYbkQ1jWGsc1eJ6jvK/4qcSKedhaQkXFDPFVl78Lt9cC6l8y
q7yBUoh2TiOnPgQBUjsxLvanvfivwpJwEXQ9j+MHbX4zV3l5wgX4t92vPOosmvoTDHhjleAXxUhu
Mlpnz3+Hym6gBcUEDgvqPleyfv+QFHBkKblcOBFZlrLwBxqq+StdPng+XO9szWHcMOz/RnDsnYuH
i105BY8ImXX3bQCzyIgyf143r2aHoVhek9nbgOnOA9SL4dj4snQReA9lx113UctaGjBNaiNEHRlN
EYQBGdahfsG6Do5uWPrR+86qFzej6/DJ6zK16w1am+5IB+zybr+LGM4AAPHn648UPX3o+MrFJh5X
4LXtEpdLg2cuJaN7A8N3W6eBDQ4BKQzpguNx4nNA4rgju6OddSitVBl8Npj24TeGXSAFIaeIlTas
dwLJSBc0Y8tssyhafy2bkCEliWnALtMcqy6j+Mk6lU+t1xAfkF+Nbs9YvAix8Z7gmtMnifsOc27L
Fk3NBUvZS++L/2baEzGyb+6YCaT/b+feA3yBa4L5+/mFJjonqFlPf4wIw/2cQHGCPlryGL4EcuWT
S05WytV62YXfT3TsEVXvxnLnwlXAOu+O5T3BeQqird120+siWti8d6dRdIrrfb5vNLYC/IRuiDIO
ZNPkz+hO8Xv2UcGW7fH8Q3aH7uAWePHta2BQMwJrP8SbOncKO8CnDgrFN0lF/2D0YSBbN+PYIrpk
GViE31qkgGoGZf4Su304/SkVt4F4dc4Oyx15EHOmn+yqFh6EG5vqMw+LUnA969fb4zKuHixpluAK
w1jB+ESve+QTuOftTAjB8Nn7/cnke7eX06Ge898N1Z1+uL1Ai12Ke4dGnXQwCqF17o+bn9zy7qUn
ztUtJAUIkymYa1mDD5jyZsZn/SvKbSReaio8k6NgwVFFN7qSRKpY4TUGJHQxI/3328xsaz4e4WnZ
0gc6Y9c1sIMfIU23tQFmTCYGhjUaZdd3auIuZHMh8rP2bnyVlYpB1yeiA/12nruIVX4o4pJxDP9i
QzPKPwBLwPEuD8s1ou/6BDVjU8/a0jlqCc3/MLnZqKKyQXL1jvRrDMq3M7Ru+QbjLdlILiitw3/Y
ErqBVYvsKC1avAWF30Sko0Xdf8xpZrHgalxgrF+iZuGsrRFHfKEozI7ps2ZdROLPQaTAtaHrc3ML
d6cjBj87dMZdkSg4Ta3IIpIyt0xSvIYS+iPYNmd/bVzBxg9X+OiPfIYQUMAsdZjGXdbwPXVeiGiB
qB3cxqEMPrAzOK6++Lqiqe9bnYoPNZyZ3l4iSeZ1PNhw6YZ4lT+LWjDE6DZQB7MF0zmCpNttrOVG
w3bpAs2KO3kgaGDbf5ySraAdd0sp1Wy4/K4STtRDNL/w2ehphjps0Dxky1xtb+H/kQXZcE2o+/hq
QbXxCj2f/uOmyNkkBxtiD8Dnvgg7H8LVwCjeVrm2+y+zZWG+H+k/9tHuedSNaV70gUjMHAENIZ/f
BBM0kI1NNQkF0H85iNCXUKArW6/ZKGIpcXzih5Zl6zcJOLYoOnmlZBPTJ4PDgNRx6OByARXBt86U
cGA51grCqFrgzorKzA/PsNQ3T2hTmhaY72kzflgxSnJkpcON8+/PBhBVp+vr/8GmxWoLVj08uScX
3dHN+leIeSpVVKWIx5IAOqEESp1ErtBg2WzmwePvavIpx14P0sPa/iuV6f2fRzhrcI2dxUsNvAcj
Df7zC0xdu3YstYcwBwVfje7C4h7LR2B0ZZqTPcx1JLNkWNJyDTofqzxZDtWOtu8pBFjTNKHJKNGw
jsysDA7WIkSF6FcWrT+9zueX/spkzE441UTBAia2J5gEzVDf9q8OFGb50y3gRG0LRX31oVH5w6EF
NMVkOMy4I4lnJIACpTkeJV1zuAm/oAX07QJSjBAeHPg8PxL7Wj3jtTxZyvsPGTuiR8we6spVom7K
Th2FHQtddfkPJ0mVSQXodZxYfoiHuZ4WncXSWBeoQOfef00DqSoZO0tu6o7tz9gSQlE77DjAJg+d
2luM3ECsl97AbVeY/GYeqOscC7MNop1d5FSk/gk/unIYJHDbKy9pO+WUBcSC6ZYD3P/PCtvtD210
qozQOa1hA4tt00aodyQulKCCgbdFMVDZL4PtMkyG++lGZxQvn8vcIzowhfLjsGD74X4g82NSRfCF
KZH1fPnmduHXyNekVvM4IRtx2aOsChRYjXNueHvCyPLllNgSRUMBlk4mdMK1ycVga1FGLuAEu30G
J2s87/tkt5EBhUZeDFB457Vt4UVFXodnUuyksE/QHNruE0GNVSaAWbRFqlPbpQf7Fxb8wgK/wumj
tg9gs97KoWktoYlPyYCW9KxNZHITsUr3vC1fkZCDkbE6JBjYwyOAe2DYwiOj5F4EWCWmTtejBT28
JE1WTCYuIQgrFO4adryyDSSZ43YnYd4038k8e/dHbce21K5UfPAwnH7lwPbIyrRZEKgg+CUy1M46
5kNetyqLrG3T2NGwHrgA29tBNImVHLInxBuGDK3O0hJa8d4UyNePFFcmqhY/nhSJXDx6aRXNZclZ
UH8eAzc1Kv2S3wWp06uCYjjF1xrQUhr36cBJ90ybSdktOOLvn+O1JnYhLhAr2FGpazkDSYUIJktn
37/UXXlf2Bx9yH1ZAAdJExmHvIAXlIvE6ukPfSPQXNLFJ8YZ1TTibdUe4wm0LQre1J3TVVMkvDnY
+q6bacWp9Cqwp9DseAf3Jk/VUJZRebEF9MeQPFV9qw4c51EF4mM/9l6VDDmoi3uUfe49ReKWKErs
U0I7+ctvKBgWtXe4VdKYatmRlZ1z3NLWjBFaNZZBELgmBTlssCZ5wlmZ2JQlz7oOmYYYvAbSTo+9
0b1/AnauYtTy2UFc+nYjaLPVfFdWY/S1mlEVXRUWCnWejzcGf/QehXWQEjAgecR++YR/C3/Zmz82
n7hyyJC0xjhwKYP7Ace6aJWsP4d5pG9BMw22Nrsl3sFpwTn9Pi0Sc1kkagVpYJiOE8Qs+mVSSWBM
RlS7qE2aawdmF5ZwCm9oTA8LX/CHu1H+UFC2E28nlyLurwHejEmtpBur90AQxn/qCcUXD/VKwNH7
HIWt8mKyWispeQ7AIHuMt5VC0uzXwihMEXTtR43FnfbuCk94Cjw756+3OMAWDw83wEMTZP9zCPyO
Yat8InIYTuxrQTQWTkQZkRzPP7VWXSe0RSlTq/hwhSZSnJUN6qM+uRCe23LjQuR4pvX9B4hevq/8
8m/LNnPCI9TQX0tJ1B8it3NLz9MFOLyhm/zjyziOByvEVydNNbbza7aIvoqYNSyAUMLLvAaYgoUj
bP4du1vZ3reAIzjWSR/HtHdt+xG3JxC82qWxq9NYP6oKfzS7/zbbbI7azyV/Z6AZWagAn2X6/A+h
mKRn7xnLBspRlXW2WoUSz78RX0FsFgW+Xvw96b/r7UJLcqg0j/7t0OXALQzZy/nS0abUhPkNwAUI
AEPbmktw/XedclWSPHKxF103OE8BGJyY5lIF2Y5BmM9Tak28B8Nsd7xr8Z6M2pL8WcoHnbG7Cz0W
IB9k6lk12Dsr3xJO9fxgRYrWMsd1xdKjeeTxfU0XauMwbKvsCQJ/5q49bqv2HizZSMJYFOLbnbdI
eAA0b47B4Jc9WOTSJlIIX6UVIFKHqGU2i6ECXwvu+yVOvAHG6aNyLZpbbhX5cSyKVEoRn83F7NIJ
ijDifMMxWkuuoploEtap/J9d3ZYmCd9rdEDVyuREMSGbjUMNn8l16xaLayKLg7og02kVmGiFFeyq
WPppt9t8VJubvCAScifI6nYwyPWVzepEw2lcci6/Y3Q6cfPYI2OeJbsGvCu62REzU1Sq+iulLz4p
ikVZRrh3OECApOaeNOR9Zi/QR0PLIA266HXVkXk4Pp/AzKRUtVxQQLfSyfol9pLN14oYB6CQd1Bn
KjRIzfisQxpRlTKWBDEcVcjhxfOHn4aAOYMKkgzGAAOgDr1MxLVXfrTLtAgjbPF/gJuE5uYJWHYk
Pv1jiBgiA2i69ZeKEziY9ce4A7MM1tjcJIql7eL+dYyInoSvNc+mFw1/4J3wlbVxeen9Das2UDBy
vGNWkzNTk39hgRRKtPn7hC8m2bFha6pfX0TvjEtJJnlUtVjBE/Z1aTSYfhSez9SF2s4RpWSBNP5P
SLnzpOQiu6+4yRtN4uTlzDokSMG/VI5hKqD4SrzQwD9L+opin70DR+uHUXT4GVFAs6r4kfzHmS8A
uPN85A3u37p6dxy4A+LgbLnLDiW8oukHMt3Og5Qv2jjFB7udpWpd4raGDd/s2ecm11KDnqyLPXqn
URsMrR76dxJxhgjMNzbHbLsVebkn666wDKPuHfwkNEY7DOtFgAINZjMCUSvmG/98q+zp4EwrdkC1
EBcXecPM6AWtxoaHMwKX3qAVWbbVcVzfKvumiN348rPVB1rY3h7DbEiaHBGC0dZPRxTmVjdHUEK7
rcE2bvctA1NPWaqRqlPva7uEm9OgXt2TdfW7KBod03tk8zbFBa3WOZtxoux5pBSEaDp5nxbPlmd/
wvnyOOlD7C8xI9PQ83ZrJ+cmIJACkIWkbyZW/KaArOI/FYg84wbdEXFQI/KuuvoI89SjFY9jBjli
yTL2oCkWEnAdcA/uRmLlJi8DlticWDmV3JYXEZDYMrgCwHUcCdt56BLmGrzSZ4hIsfIcbJjGFpCg
FA5UYpr8WQQRjsS45uEr6nHlxXHkLIE6mpgjroa/l2/6irmPuskIJdGiGR2jkz7b/lbXm6kxQ1ib
4kYR2oDG4Xb3R2naphwESPyJ5YXs1UtUwQrlVNceh+CBlhegzvXUSWjmQ0/p6CpifzfAFp69Pn7S
4930m5lhAvgOy33D5YaiFoI4OzRl18IxiFJqEwUlrgoyel4lD5ayu1GbGzcKsoBymaI7MRpVP5bm
NoMQGh2wiDNlxb1W61LiuPJ2ZEibD0rSSj8BXGktlSDRd2cWOe1d/un+uKIB2NyxIO9fs+CLtkQl
z8eEl5raKOiScq0uzudneLPWfHoXaNe8K1O8QYeU/VN/SEoa/5zlwcekf9PlLJQL6n70n36GMAGo
tA5lBoEm2kOwOnWeV08mduW7332riSIOcFX2OS3Ph2nhkp/3Xyq0YyqzUiZ6VhjcXp6sqMnYwuuv
m+xXwskQlwF4HWVhLwv8UDMJtT0fnBR6bgOZOVNcfFgwCPqZGbWcEUevWTSaGSRSWcCpvXR8SIQD
3pr6c6t94BHXJs6ORiovfNuMFMOR4h2s410YPJ7i7YvTQtQ0BHeHtPXS0WxfGKnfVaKDswcp7me8
JWHlLpcaFMSkWm2VmtCe18huUimRCn5lHIG5RnVB/jz7oKlDo8raYdfAzronJnkRURX1/OQYsGes
m4QVZuEwL5ESI1VIexBlrvJjA4jqaUNtd2RoXP/JHe3aBF7PkoKQcjMHO5Mj5sj4Ga8XlE2EiLIr
PvA7njuAn/mqgBwrT9DXtIhyTUVv6TyjLQ5+zuwbu51XpS4mMLOpkvep1dTMlSjtAE4eVt2H2mtM
fs3eMeS+6gY4PvjYKq9S9UVSCzzIr+nia6FgcH+HdhQNLvM+ovGTmAYO+8y8hH0Ut0/pw0TqkrRF
P9eYArzpxMLQ2OgSsZN0tuvTSuwDSya56gSshvMtcjlu6WWzLLbn9utln7Kayu3uRPzbDtmPf90z
orDdDGySkSuz1BX8gCrxnvgNO+SSB+myO5usuZywOmGVnGG8dkBe1q5VBlU3K+4x3q9TrByCx6v2
JLlRqux2Js2Wc6BFUUUJdj5zyN4sT85jpxY2MRcd/Z9LdNMT09SLHX1egG2LC2BZx1GjN5Ib62j4
h2Qc2m1N7jhdo2FS99IOCzUMY6nZwJL6voffwZlK3oBOAPvLgxMGaYq8mDJn3o4CJ5HouzvxWU0O
kn+pTgpnFCYFwnzcDsAsCNKz7mgJLcDk5oCCaDfuQ8rziNqmXclUpixJ77GrMMDBFxp/quL1sgGO
4pxyG+CYbWiiG8zPprwLC2yPUeHXUBUfY5XQ7ic37eghJFvx4+rPnY9iNuls6Ac/sdiu/fbgNuY+
t9Kbq9QPRKWVeSkgRKkR2ZidZFL4VMvsyVXjLKMXOOURLqTNcIVSf7Cqlg7QHpnRj39M3PR/Ml+J
29aVoeXPfpanYL5l7oQZ4Yk1RyL1ettgtudeZrUpacavGe8Fwr8rktQkDrlvphLhsb86effyMFgY
Zhc84QyDotv7juXJiYgQEHLWD8Tu9iYQZGq3zR/Ond33GSrQoFzDU76xp4Pp8su44glFf+8bdHYf
rstBfNKggDQBiMySVKxo6YdGGV8csO7dfJ+qt7sDVMdOz2rOYTemI3pNUTT74gcZK+f3xUy8ShF6
BKw8Q7SFa2mynW8BbcUWZdtfxSi9oQ+ZO2abvdB2azzDzy0R4cXdLCCDR8I83smh+Se9fDd7kHto
UxnVGwVVUxP4rXBXhY2EKGUv9dtj9DOf7xl003Za9pnQ6+nzaan1qnc+U0a9NUPQ2S9ayDz63kdo
Gefdee/fOi7iaDUAvpKQcK8YYGawU0QEFsYyT122l7krlyzdBhyeUROAi03qt4EmxbfAqLxszOEX
LvsaBw8E/MCucRe6Z/2KVUag7VMCcRGTpe9wPt5vocB6G/JwITg7tHY0RUmiZLzM4fxUsaxZFLUi
OwNTi7pC861FMlbt3J82JnHkkuGbvaO6txFsyge67GUgaJRSAYj0YlzBs8UUNe6D4rtNnRclFmLm
2r8dPLOtBkcdfDe+I4RuM+3i6fMLD6GYdmUgtZVN6UEBLdGsKLTmvhrZbuTPjqumz2v3nD5DXGrD
PQyptT1SALL8pzr+4MNJYfkTWfuZUvoJ1yS02VvtsYHptbzXxVO7bqEWwjgm9f+7Sis25OSK7z7R
BemUwlF8yuTijQsct9Zl930D/SYzNkivL5GtuFlzDWCwuokumrjRjpPe+81J1y50oKFjojtDA+wh
Ld8VThJ0VVQ3bS5SxiRDrr4StgvVsXV49M9FGDOoEoQK/a+frSpGB7PCFYywc28+8OUwIHnRU0A/
fCzmLZQ+GavutS6kDwfq47thkOHfPS9be6OuX8RN0LnJKTzznMIOIsh7+N5S8xM1XlyH1+xL48fr
ni+zV/ZCA86FUSDjZDOIdnqJTcntVlNNKWFtwt0SClfsdxshk1IEiEyaNn9fZ2/Q1352vvKK/jnz
4YAeaJ7EWZV5ZZebK4klSf6cP8iV3N8o7MXxKfG7lB2rQNf3oSTe0p5pG7uLghzCdCfScNINtl/u
5Bq2dRqbUqMusWpoBzOGPFEJL28e6m43H4QaMI2dhXppPEWQjrwbc+G6XCjfMUo/8a0ISB0/+oSd
c0JajE6AHF+hDHuWlcFQCyzxv6cYzSSuqmswnUxe4pbyemGydPB0YVyMvTSZaKDYdZt435n56tbJ
04NFwBpd/0TFvlzJf5oFnsOPZmyrdr97FvdcNPb/pV5e/5sdR3FL0G26c8qcWqQdp/vB6kbaNPqV
OdfIh2BTZg5PJwTAJJaqQBVAzYePFJVxOk18aYwP92eejyWpkbMFFIdoFs7PeQSPs+wi4bhJN2v1
YrBVtm2WfsYkgdk3cTTAALpzmVLIjYsaFfDEA8Kbr0lMYzkryyMaUU/ccu7QDWBT6rpfymXxKVgc
OPAuYmDAwBJ0hzTZ9f8tIciDU6tNKtcP20QCTpQT3YOaL8Q8v3Ps3DyCCucGZC1LcKoJsZDk2IdF
nsPW8engBzB5/WLrD+3mJ7gTVe91E/yHwk2MirxxLrPyOr+R9/woDPgbA/R6i4MINc3zNa+3a/Uo
iWyz43lr2JN1wWLc7c+DrP+dGbvf3WtevZNXApa4O5cLXiU9jVBTS5/V8Zhicb378+aiABoEPxMa
LQ6Ysef95z3Xwb/M4NzCkwBqMtM7lXUTAikntsXSGso2WufqxBnfX/1Fv5NfUjHE+H4phnOa3jcE
X6U0MSbKTrkfgP0X3vgxBjiiFN2x79/VojmKuLj+c1iuqECeouSUTKefLYeMD9Q/r0MW4tLe6qlA
ElQmxmGCgUZzlQuuT/iWgtx/ZFb8jMGrvV2L2dbRFB3To/hBSu9R+HrrMQkVjtDiFAjKJjh1ApoE
Dv0gMEIJOjmoKzf+7YYJD//zq3Jph1M3FrNHSQhohhUsQHRwpDf1s91hgLsK9m7s0SW9i2VnUAzt
2BlzH9lunITB1g9I1zziM/N4YOnd7YL7ExQilGuNmHjxDVfWK7JN0IyAi2iDLGLqgYBS6x3W2Vgb
OXFgWNWVmnsucHta2QDi5tjRUHE4LXC0lod8hfnETTO6cjNho6XSseinNue21dI+du4SdoOt5vbP
3hZmSZ3MH3jD39K1TTkMWNrd6XMNbUhDwmGzfYPoGUnUEzxObzLqhgYgYfPUc/Fb58MSvLOHxr5r
3gDcNMORA6kk1SCilU/JWG371jgBbptWJe8CiLEulwAqwQxjmeervuaxLn78y0CxPLifYaI/agF3
vKM7Zj5FlHia6CmhTd/Zx8mAIZEcAO00AU9JcSLx4ggrtyOmP0P3SEC9qHCX/CIpSmBwH3elUcCH
nU9ypOoHPm2eW66l14Hyv3Stq1tpSPMoevMZw2M5BCOPfLdMy/EWr2HulCSPTGY7v2DsYHp7d1/Q
AigCTCsSMwbGv8LjuXxUZ5WQbLIK4VAWSsUyLAj92Aki1JAgsdIe7u6PX0MZXQkwck6y46VGweO1
B2Eqz21CRuV/EXmE+HGcxQK0i7u2ZkZD89MBpiVU8hBZlEqD4dPHGWuqto7KOFKOn6lCcyd7Miul
dvhlF3Uni+vG4pDH8ypI97YuSs60mUZ2EW5Y8IyJ3Acs4qONbmj1DaEIZg+N5pPkqFRRNsno1QUj
IoxKcEs49H99jKwLM1RZoQCP+n33Qu5FcQSO00qf+wT/j+zkm2n9z72xq/pqqe8gMt88If2mPqkp
VZS4rz5xJz6usTlqTABktwdBnboURuiTotN8aGxEB7FSK/+aUOvzXRhPp0nXEiwjk/HtbADdCtyu
fZNOTkUzKw0K86pyrsdxJ+m1uH60gi72G4y0Hyk9QarfXICbDgG5KkPLfsySquMGUvfMJ//43op9
MrGGV8iVX4gKMeE6LAsd2tSw7OZKphi1PnmP85qH+/q9wqsAwEgMb94d+tWph1GWQQ4f5V9BMvq8
lk6enN6Q4VxEKtojyDl4d+EBVoJHxCXQb7Eh5P+LeDCWKFGiQj5k/ogScqbSUbz7Mk3ppokny1i0
fOnEszQZmaVkw8MTqIzUzXejmeA56eV4bZY+sYTH74CSQKN5ydIAEU4lULDlB3ywHZ19VGQQfq9T
luHqK77WzVY75wNpn4D+FkdIleGLJwYkKSH2jFAaQJpMcTNFciLVpX0ay8aKuF++MIeetvrnYg3I
u17qCxNLXP5QN2rhFF8W6sxiURCq4UaUinygWYw8iX4eftMbX5gTQF7rB4vy8e/NMvtasmEynaL0
mOXGwWHG20bqfRKxjMRRRFPn2TdHDFDVIXJCtrsLid7HhQu3RB6Lp40pBmrlAARD1dXTxsXYknKj
qs1++ux7Hg3Ze6ymlidumfGMoUs5JuxqoZzS1z+1XzOJRLYqFBkIMf7JHegvHhRWu8Dab32aRaze
/zK8C/M358TKnvCdorH+t3SGSAdq1MpeE+FRM1aCqtAO9zpaF9ZLy4KBqMmcGzVPhnpCozh7oYwP
PZ7fGN8GamMqZtOFJqR49mswlN0/GWgDAVFB+o4c714FjzjxXBrvYEs+tOEwMjI19oHqq7T+PAcy
IGPEwOsA1XnckZB0hrzdQYdnallDT3IPr2CtwbaBL+Je/C8NULKQQuPSlmVKe1QROpk5sZpYvlGc
EJ9QnFEJfPEUFW14EtG9GpEI0cJeH+yhFZUc1GVtPh7d2OCDlmEVWamPAS2WlAYPEzJoTKSMu7G7
wCZ/iYAfkLoruylLKAr6QESh4s7KMnE687v7FW+Rs6fxOhWFBnagnH4yric1LnuxMB3co0D3rKfz
DlhUs0WwXmrP6c9gFF08t+e6HeBBYMZWG2k26e2WrHkIjEyxKBcYBoPJbdaFzZqERgXkekV+J37z
uxtBuqXih183ArXXMmGwvHy3w7zQAoktsxRqBmktaQ7RuYFcTTZWevG4wy8hhvzvPncSIWyhpERV
VvX0jAnaIRzPnYl5hlachKOW0vB0kESRRzyCL4u9fJ+VqMMHCmCm73sVrAPoGEpMOV/mO2JjTISV
2DvbSeIS5E1mL2+o7hciNMK5zDDQ5lVp+yipuz8yEDXDg7mE5hRtVjhsbPBPRwMVP38KzYaI+dn6
HeKgWhUltYUkSXspju80bj7pu/vzNN34VFTtMP95LbC+KTYKU1cGBQ9AymK6bIarf630Oi5AFbXH
dCnxABS39ciO+nLgYYFKMBhploqiZ9MwpdFwKqFpOEDFJnBJzehNy3n6biRifnctqIRr3xRoETDJ
tBhfahT2beA8TWXI6NR9SmYckzyUa28UVYVDQQUD5/8CzyOh+aKuFDIXBb5O5x8Nh5BhQcJuXWgj
9IH4PZ31h7Wf7ur63SaxEi7+aY15ipNWfDsVidu51z9n/LpWZWqMhnkhQxP6EXjb8q4fUyaR3rKy
HpXmVuDY1VipI2KqZseFVxl9K1oX1ZU1fCBo7Bhb9iYTbdR/+N4Bb0WWO3g2v7oF2zX5ZTHqVyr0
ufX8d+tTlhgyiMCUf/jQcqKUW828R9UI+R9bAbDGAfIIwoy/gCBv3XMG7ENT9M8P25+4mEYybuxk
tk48T3JFFqGqpJ094AhpnVVPfOCr3UjeuB4us5OJ1+XWQEROkdx4WnWtyjqREjoBFg9osMN5yzW8
2duwiyYZIIN5GIJme0ByPWbybIuoxa7j3sEJ4dZ6rZJ+teUGcunzX60hLUnWq84sNC0U5GUU10ss
yHM3h9B3HzMRIsVg2otb48em+A1OHN++2FF4HG+zsMXAvE04+FaZUfDjPHhQ3x/SxxXw+oysdb9N
bcmcpu4MoIF1qFcw6hmBRX2jpoZ0bb5ftbF6r6Xi6A94c7I4ejIFJLQI2qUYhud7y/J2Y1QaMkM9
Dz/Sb/0ZcVm1UmSCYXhdxnV4l8tiWZxKrK3fi10yXwI8CqfwSYhiWh1QnOrfStojavj73P3Kgykg
NAdbp0BCeJIx/ymt4kFrd7zLwwOarvSCPVm4yGCv3sdl9ZSUF8039iGZryKvVxFjq2dZ+116ggZ3
qwUeBk1dx3sX10ySeyNKHQQe7zMF2p8QOQvUMuYqlxqFT/ULL/Ofyy2K/GQZ9IkgZaXLvwvNbXH6
xdRtMmkJy3efvMgi0R+DtlM8bCRY4x9r5g2k5Xu7cQRx08Ui68JllRXtQTzjSbQqm/YeBdxZnk/A
oY8seLwRNWCqemfYgZBgmKyjGGKOzwHjVK+6w6Skww4+bR44eFGBJPSCU2xs3AmlfV4GuCS4RB3E
om2lYqkfxQZizMFS+gbOIm3RM73eosdp+p3j5oxbcRPGBJC308oIZJ/a1ePTyTuMBLc7LKzAZ0EM
+dB4A1h2idqxE3E5e+8RO5T+r+ZkVK/7OvK2UGnxrGpUo/TS0ena0nnEKyolEvMaddcxx1B65/Rs
SfeNL5DLiAo6Akig8HLK5KV+z5Xxeulzq08v7wQPBsR2YBdwQ7n+xWf9AbwSjaj9F3UhZdsBNwXl
QiD651eIkeMX0I5Tjel0ZOlM9hrpzclhZqXSgnKBX4GOPFHQsT/o2Rc8ygjjKlYfAIngHShHCe+p
insNx0tSuwZWxcV66CWVmDUASL7NZWSKzfX770Ee5Ctn2w3uQjs3WZk6fxs3J0LbzuYaYHnPITUB
pVzage9OTpR+JNxDFM87rBGZe6vyL5laehM7to3Fz9SWvBNjbvM43SxGr+iktMjkTNe67mM7GInb
oM7Qo8oRNsCO0dHcPwKxg3GZvPrR9e9NIdB5YO4hQw2O+LQGUWEZMFc3gBKDXzBBs10KWfRSOBFU
gHLwu22ciJj3CAbkdmSDAXCganPzRQi/Nchg0aOfd03UPyy7h4mdLvu1a5l1ENbGf/czOQ1e8Bwa
KmOrH307M/sMnZB4ANJ82hi8z1oHoxXg7UwSs2IyVpmD3NFQnLJqZeLH9VSjuDphI2Lhlx5C7jAj
fdpXjmw31jiiGmfsAX5J+S8xYqCayyh67m4N/E/qNix41fdGjk9THz+eYeZRxmi1AYVF30ZqBWuM
AMC9pLPocLoeJsTFT1xNa4twFKwBqcMPfyFG/pDFujqpAiBRNNXp/XPLtR4RZxiObPues4/Tz+KD
UrX+++5vWTJrbbOC39Vsh+efdKA/WxtGnzvyj2sfFl0sgZSlBA9ZUwzvA3g9t2KkEjJzA1QTNvj9
9hFVqJDkC73O6iG5xqUkm5ifV9rb1oCrFe/KYBYPunM8UiiVLSxAco2/E5rUT2gn2U+utvuHvqDL
pB8UuExazEUJ3UCRusZophyh0Gz1BRhpVWagAn8xbBQf0zrp8oXptIVDQEY47ByDr/GkikQtNRRs
AXPOQepSfZfI6G/30od/+zvDPvmdstNGNcYOlwTEH+EVlh7Ez+VkSV3uN4Wt1+ndZ8m2xcb0u0RH
PmVLn+88eVI9ylGOrdVAjCQLfHaPsbiPN6bKgEVKU9mzyrJThZhfp4+0v2h1ob5T7fB8+pSSr1Eh
OBGcLKmQFxOxPsd4tx/Wby8H7sm2Z7ef3KA3onRqacsELHMWMpGYgHfCJ/LdoktDXITzVxUIogoI
cW3nyhuOE8bDi6OvvM2nv64xeJaFaQbCECsfwJSpWYZwX4WtENqwlU9H4LM4AYHS3Ataoh0wfoot
bgMjsSs/1ACxnfAKMvRetVTDKSsrVaV/0fvMbb0SdvrhXurkjZp92BVr/RQ9RtrNIdUI1amGU3Ka
nUyUPNOihmctyNBUhdqxKTKZKP8qNen7T4Pfurx8zk9ZqtJEnXTJgIxbR2dojaR6DwK81p/nHA82
dntgDBhI0c6ikpKXqCX+00sj7Y1BWSwywUGCCrDL/a3svZYuo2ZeQgpePvYYoMY51sAVJWnEES2R
/fidF+nRu+sDAYZxmhFpfkAYzxTrCeYeSS6ftM7l50+gtK5D/qt/IiURcWjAoLFOe+nV2d/qSz6S
cTWiHGK1dQsqwaLwky+lyQpEU2/F/a6tw3gb65rAVHUCZN51ezTeiwXzo3NgwEih8Co9o5ubQsO8
rJkvc6bV0kz6OGZlD9bOG6E9TkH/ira2g8p/F/TQOw18GS24H5cp5/S9StKi6wMm2RL2xI9LVm1M
8Q2i71EkzUUW/XDq7vlqKmZD4hA4ijDPi/w5bFmRs/zagNEcyy/IKXJKfFNZy1BJ3o5h4MCewzWO
4O8gdqfYIyoqLyl9upGqf9qe5PGelrTEa6nOhf5uDt9kFF31xOhbSJozEUBrKCMmdjNOi3s3sc8r
0XT5YWdhQYX9MsEKD3JvQRr2Ruj55P+DfzfWpSV0//A3KUIgKNuxdmMYts+C9LuI0JfK9kz7Sq3N
s2e9XDcdrNBwWAKvyctjyy+qoFsPiZX+x3k55kHBbiBrsFa+nof1f2YLJkf5DY8IU9RzHSLfiBi8
WSkcH7WTtCGO0uVa5An6Z935Q2ch69AiRKAQBZkJP4DlJefvT2fjvOrcUnkN3JntV0oRYcBapj5o
R6a3hG4Q+IRPIqcaWjsU/W6zZk/QO8+wwtLYHBDL16XucAkNLZTAXKKXeuGee637k6nPjWOpxMOA
W2bPXqpg8GEKixprBBiBQxsQd8km3gYHYZ+w1UA/o/23BxFXE9TESEU5X7kqyVlm5B8OtGOPa/HJ
YO3JZaYI6FwyyniykGuTUiRya2npkkMgxzSzFfGFB3+oQevS2vyZHbFIrAOI1OmLGOo9396keKHz
Hyt7jMskCr8jFMHYWkpDs9vz+4Bjb+zDzuFL4Nq2TZuE58MaYzunmsb+qj1nIMceoEVMvKMXNMQU
k+nzPDhVO7kUh94+PB03+wj2rO/uGU84dBcW/Th9C1jHBM/7pzxRHzCG/bvswxCehj+X7s5ODBmq
Ksr64REHUDZvT/Z3ylUnZZ7j++HehXPufmlNdNVvpRYfFFIXtRJTX0Nu32QEPBhHpjh0P67kLWN9
p0MMnmCcdpqdX9uZ9O7EUQVtfzYYBCN+kM9Bmew4hUV8LJHSxPxRZdc40GouPtzG9Ii9DQzfrgn8
C2Bn7D+uyx56103fbQrrYXJztmZSFLFOYnFwBF5MnbgFZJ4pz3yhzEgqUug3wVFfAQTvvKT/JW4l
GkG5F6NULuocj3M3A8+ZyPvGkqVJH4j3GUZAc1YYsKH5mHDxeEz3BuPu0bsmYp4WCJ6Ua+fWWgo4
hvId5fS9CsRYZEadYVfyvAwBQ3MhgXso0lg+vlkeDVXw1EAY5NivpfCQ/6gwVhCLK1LsOdLPBUm/
QnHKFhcLNv+4lliNPMDDo6xzIHUe05H6V7YfVB5TRhJMIxB4oe5iF0GFmKsN7/rUJKTl4BDDPfNi
ygjY8byMm7njthcKfpD2QVrgxDC6mQyDIpbXttvvKV3aA+nXMRRq7vXn0zb4SSM4RKUXz38WvRc1
0JEiufA3QorslAo3cpNM2dc70UbKiytnnnVYgwloGiey4r1CunOuXFB9bP4Dr2K/v9G0Ip8BbNMh
mz13rzGKSCd4gpqUAUCqBNZfmUdJWIWfg0B3YXuIm8QDQ9uyRiirB09mxgk3Pa5oJ/88cgqfxGUA
kDM1Xwq4FD/T/tJoZoDQ5mEGue0LGviEygc9gs4rbqsArjnsY6PoNV17ozTroluqeVsDdebC3FY/
O0nd3x80WpD29Xb76EPvO2RP3tbvYWNqAXAkHryDRvOGQhoqoxn5WB0n812NpXGysj9H1Z0oJ7Q/
gZXSxYPR66sOihfYzHewO0o3ae/GaQjdbTPTXFCMaZcubPRk79dD6vimZ7IKnZSNqJfbmoyFfdpf
nDoMGcnsodef+cp4bDCNb07489KId7BjEEfHu697pCKFdydGo03La7ncpg5zruelxSGreHGYkZ7l
u8r8xuMeNJTrkxZAovL6rD8ChNpY1zEVYAVE59BflkRAUexS3cfb7pW/PLDxbELuzATEgoTC09FF
seKbhiMotmDbF+OL7Avum4P1xZQbV23NwKm17/euUdgqxr+1kVZs8SYrEy8xjJQ2ctMF0zI7/Ztc
gLCZuwtbBlo05ThDaZvKa6wAW+oZv3Ns1CndelvKjjDQkYPc1SzedhEWVd/hv9yTDe9+yojyn1Nh
NIffPkVzTargju067ZF6iyqZu+8EZ93jTy+KsSWSIYAuTgyFuors2CHI+Dabn0KosjVxZHM/6gSR
nySRD0ABi5VQgHmiVcQTqszykoiZiZ0Aep5q+2ldAymtaBSeLuVhApOi/772GmSBHH/GAm7RrmBp
owNj0ToTHmqTyWCIRGovfd8/WOOXlbjlzrrzohom0DlZsKiot895Zc8aCz6BMfsfnv588Ifg9Ghd
y0zY6+TqKO7Y0ES41liJFOryITG+ZBUYjOzIx6/Z0s3iZhk4yAYpLErKC/csXQDATQeKMqif0luW
unvIKbJlr1LCqL3HNktWKyqT0Ux22fDD0FJc1i6MTRBhXAfDqyGROG1NwG8wCLn/0m713FE8S0ow
Qt4cGPtBqULhK/E4TVV2niPMfVqSwQ/7jzxgcmM/Mdj+rLD3OP0ZrYEJkD+BbiSO8S5yAgnkhjRx
/uxEaDaxaD87gTodRxMv+KMQsWo0mAFcpw1DfY/iUAydomqF/XZwku1T2Z0Hkud4+3oSU/CGUoAg
7KKdha1XSapwP4BnoBTaC8B/sKSFS1GijVDaWvm/Ux77aUSHSs/M9fB9CRJNeq6adS7SFeUeE1+d
XB6P9q95h6JGlSD3qsu8pr8mCufI0xeagCpQX4sdSNkfU5b/DeQebUE3QJxMjHvkqWJRbMGSQ/Kp
J7RK8xpBq+4ji8qi73572tjILMvo8hzuZnsjama2QZ9YubQ+nVzcsfn3JbrplEq9gZZuIZPFNhXC
eG7rg5cdpxUkaXS8Ot5NGvhETxRmIkL5oQ0+4AjMqyOvDVUF63C1ACrFz7LpVzLuosPdHor5Q1iS
zqiZjYmmWjgvPkW2RZ7ubk/BF/wFP8YdSMIZzMZWZu0nhmB5wAw0AgddhCZmojkC004BBLaNK1DN
pQJCAyrASUhP7ogVEa4UCoDl6Paf9T7nC6UpS2c9e3to/rl+p6eJB+4XC8830KU0ak4IRBQha/Pc
zDE/YP8imW2KcPyJdkY+GN51Wua28ywFSCEoqdYJRoxMLdqaW/i3T8oJgiR7ImbXHIt4Bg6UzO99
fS5fxaWhxtNaexgNFFTMyXesWBduRhD4EStT6yqGCa78J5LJt6Px6mkE4wJ9yt483baSkYIkQU36
mmg2R3PRoVeRZtyYXEAuyKKAX5cE9ZE/6dUpP70V38Ney86gG8CoMRbSmsh+qKfz6gf4yMcuqdOH
Ml5ofGpFsrBnhg9nrdZJiTzGZwN7QIUnwev2YEl2MIX+rT+jXG2/CHD6ggYIwVH6uz3fTXqXpBbi
3AOEaqov5PDn1DNdG9nRM5TrQGUCuKYUs8zY54g/A29o23yRcOvKYPYyHTCyXlxChiJ+yk2fLciI
IjhacubFRZyIA5BtbllbqBM3U6Pgg+8DlAO3UsPyuUPAH//4OAhFqW5AUvzY++c4a5ZCGTtORq1Z
nU4/7vTiviRt+K6UAsayCrPAVmvj9u1SX31ODE9sk2hwfepT3H9sPP+dOwlBQ/O6kiHZ0x1SdLUm
NxtFXizGR2wFAmdQqs7Y44U+qJKyhhV0ZkqCwNIxEIKdcLRmoRwbcWIs5mH+iFPjt/wa6SaX710T
eWSSCri4TNxbAbArnQqmgvlOHRIfBPvbYQIThlmm4kRsGPQ/LjvILxThYDw60stR54o/9bgamrmD
IzQ7T03Knvwlky657vo889uB/PgBWSZ2Zyt9HJSWYhV34cDRB0D491Cnt+Jil733CZU8nyVjwjUQ
fDzc9ib1zJqBKGIRMAgJ8m8/M6iiobGlez5VCipS/jAmaexJq1xdDrBXKRHdTrlR14ltuqBhB3Wx
D+w6Go4L8Wo4iKIdfTA5MYTNOtfmcGvVcsWHTW99SizO81Kdl6CjZgA9ilTb+nYxnnVL/MfwylJW
dWUc880xVOA9OPHVbP/3StOR8ECkpmziw4EzGZVDOQo+90pJEWj9bkVbbmODnX+uAZCrEDiU5bl8
vpSF2JojgJibDXeI2I7Z93X5hjicN35T9XcUYlOQgswQm7X3Whq3mgKQXD2XoCT8ysQZUlIXasDg
AXMhWaB6GPzZaZSq0+hZ23OEoZqdKpQdqt54RrjoYD7fr3sKSf3INaL2sttzKXRDwDl9+AYljjn0
pChLVt20T+dy0R/jZgFH4Tmt/CzHNFBcZQOKOdL9i37LgR9Mlzdu+nt1Srv66ELBtkV/5PLYdKvy
iA+AXY/9GExHyXjeW2Xru1SnD+OEiOGui1P4JTI2Fz2BpAtyfcYBfkvKkkGmf6AYK/C3h7GEe5bH
sDKl4bg2amW77y+mO7Jr7iDj5wWnq99FFbRYbGPDz12MVQ3icCtOfZRTVDUoYZ6Jdnx+W8wOU77o
nnu4ZPSRYg/4olIq6O1vFDAN0lqv8gaUWZyCMyaKnALvFHq5yFQw0zduKd9OCXoWb0UdiTs2wP4i
VyAca0Aa6pGvg4Rtm0jy2GzCdUFqtitxy8P60frPb5jINYTYtYo6pe77WrLWIvehaIe44K/bged2
26tIi63ESZ50IkDWAUsiLsYJDJA2EF85qerPv6YOi615SlcRoEdiow9JSMAyI1QN+nxEtNrB3UrZ
09y+v4FRAAS+aYeUCJa/O9yIFA7Id940mhka/i8/Bz+VjmqcK5wWDxypelx8FpT2WBOKh2EV6Lex
JXrh9LXoeS1luO6iIERFh63qbi4jqBdbINfXNyZMZxVKB2y0c8oBueomMjpPeGNP9ONioZzksbko
2jSUHs2JoMdxEDijSd3XQJOR1mlMCfubfWDN0sDA1chgQpiBhLCxVvm1wffJaaB3ePrFpCAB0N+E
j3pYbZqgj8HdhZ7mP37DxWuX5mA5XaMDBt7u9RPnhuzkv4/omjctPHDQFPVEXni/6j3dJxgHYU4L
eSdjYEACyHhT4n1AgSsYhhIlEt7biqqC16bhG5+1xHjsTRulDGbA2Yfmc9ayA7L8KNx4OjfNdoet
UNTf66vu6Fd/FGpg4FAy8kfH9gWawYHLzyBQdYqU5+V2CBM4W4Fxdt1QTyGyGFF2fOM0Dxh53ks5
iGia4vGvn4Jkcd/rMh/8v92lPv/vVPErI9zAs/2B29KSDi+7aBVJ+xbz5cXeq+Y5Os42oFz5H/7F
JHGoCE6uwzHFpuyJyuSJwj/dVCtL7t51TlGCFoDCy1GdeJIf12mZZ9fMtFlIGFZo2qrmeVxtZR4G
xgOFp7kHjY/8gc/dnhQEGAIzvfSCLKoIPmNTQcJYB8yCYQndy6VUpcV9iW0RIbJt7mtzIvmmTF5C
EGzOWO2iW3kgRWH7UMknGDrf8S+Mhxro/W1nOPvE32xQRAMi3Lk4J0SGxgGQZYhZQ9o8Krv5v9cr
MYZAx36BqfRBcf8ERZ6Ykc7QoZCM2bY4my+RnB9ROtW6/fGqKsoDSwTLm+Qxo6U2p0l5pJEKLCOV
NqpRRyYHN7CWyOLAAISc7PZBIO5uhbXaFA1aiX5T4tb7Hx7rnxSWHOeJ0D8QBKvOeaXhYhq84daX
QY/nfT8tb4RB/ZarzYkMiU+3lhmb68s8gaOD7nkuQOiI3RKBY+aU/ou7uH2W09Ulv77K95PT33Xu
Kt21bx7KrdIBFSofei8UoaW85sMc3VZwwwTMHQkBDdlErDNG/GzKX1kiHMZI6hxzd5ccuN+RpbFy
sxj5FUlniQReWgQxRNmru/EbwCcIwRxP5eiUnAjSrMOjrHej9FkjynDTCjEEWBtLIAkBbDTfTIdz
CVnfl77GfOOojpBRCs4JKBB6gdC4DrwaWsjMA/qRVRd8Sit7eoOo3ylH7eLp7Tr0+OVXfIK9jE9I
FM30bYI+PeFBGQOXqt8oes4DN0aiuWeu2jbVLpg1HDvOzOVcXVRLyMKcEMY36ug+UGOXiHsQGvx9
MK4ckXd5f8dof/v6l9zOQTV5k03cHaa357j+jheLT+RfMLSTXI7U9WHDeXkxJ5A01EGTtCe9n7kA
KSdHn3PqNES4CKCj7m9aSsIlsbsm7aPFyxSrY6utA2SgHZTfPizHrrthbAEqDrBmE2EZClzW5zoe
b3b3OZUbwyZnF2uLoGOmD2UFF1Uy0lv75xxHG61d8VY+twJ9Q7VdxClxHnUWVOPK4jRZOivtvCna
CBCO8ugI9DQ+YZBZU/dNnT4vSjJ6kr9K6jhFrCXJIcS+a4HaT6RpMBbOVBEZAslN9LaTbBobtAUN
FXP37natE5ssJwSoAAuGKinntTw9xDAHPo25q+aRq0IB4PsQPvg6Yfn07cNjZFF2R7pE/eZDSNUA
NQsxfAJ6Q27JsCidaAsnmzZWffyUG+mJlJ4wyhP3wIGi6/UUwHYQfKi/JmCut3TpgyOuQSpHbWBP
yNrKKbB20VuPXp2mGE94L0j4EJF+JLbrINQzNqsulsXL7HK2kpqV5uM03+eBxBWEWIPh6uNMOqG+
xhFf+s3lMmHkqQzghT652jVB+L1PFipRUJ9bnhDO41h17eVtZ47AQGp6WH582Ezy+aU/Ok13AIVz
AJYTRJUKE7Je55/nl4ne8+a3OTDB2Y62yzdVatWIuL+M1TOLU6OUOhiLaGyU7qtv933HuFoGtPmn
nHkmhjjIdVDF5kk3i1PpNnS1M5PcVON4QugYRz8sEh6rMx7A01iGe7RB7NKeDXaO4A2pXA8LUlub
Qfv2HEnmD32ESNakXvvKtYdomidSRLeASft8kEGDbCYxj8i7DbfDvF0jVqcGxtYW28aio6oEOdzH
Hs8+W5FgOoGLfyuyfOiQi0zcDrhCXMaY6eam4fwicHsCD5jzEr49kB7Mmv/Ib1anbgda6F+mZsq/
611aNfiDW2trfLGDPnYwSJd1hpDjAKPmpaNV22ktSj2V6c5n7Czf4qjvoAWSQixaTgXNZkhP4/5g
yHgBDMO5YJg+j4Fm3IGD8VA881cK7PuD30vGYgw0R3krxNjMWj29YF8pWsCSuW5e2xCx7TFBbDMJ
qWvmwVo7+u4HlKvgM9ibsJHAJ/7h1i/IQNVTToxoOyWDuwFX1y9FWIrCxYJxq38LMkGBFYYQobN0
tNb+wm3ADI41OdIKRMhXmsHDNGQK4uGH+Vqo7OULydgbm6igIOzZMKkWeFqIZiaLTbUrroH7KrKd
SbUhyjixPJt0x1ojJ6bm1Mh65tCujqGV2A==
`protect end_protected
