`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aiZZuAn46GlBcKbNyXuD6m4yqrf3AkOrRRLfbjUPUBDznTrHOmtgmDl6HP3/AbBGF44QEFIp5nXL
WQadxXjQvg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lahfFvzVhSSDZxrPSUML5yazgcVNuICUj5Lxe3X1yGsmVEqH2y2+qC1ST2KWhc2QskvKW9Z5X+EB
4IuZMKh3Zj8aMAkcpspFp/myhXPtUuFfhbO5l6o683zak5VM03Eam9S+8VmIcYLv2WlmiHb37Ydq
Gn5WuZCokhiJdsGXIRA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O9/ADCcv9uUAlM4tWGQc5kCnaNWkmBb5+KhORnvjKHc/88zHLo7MAw4RbNj0V9w2RNShPkDdAjIn
XOezoh+C1LGI3jIwYDQB1H4hBb0tIaYG9VjMJcb0I7wWM76deX+wssUNTY9E46R7e+cq5NRFLuI1
nJkfZAURb6o9V0yUb7iTJn0u+sEaAFLfRW9+Sjk5ntcQyh1JIvnq+3ZkAQAhiJ/anUY9HFtOHU4Z
vrXR+CuQFRg0Mpyy8F2E4LSpAB2dTUPphJIfl0G9jnxsR2pdCO1V24RzU88V9FZ144uuq6+R/bA4
RyTJ24x6hMxpGJCyo8hryTt4nyRVNTK98SU6pg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rq0AoEYJSXUic3Zh+ROLbMwPbo0gCwQw7M+4GWA4Jklfxy+l5/s5nYraSZmbcEHutEzq/DecbymB
OvJhG/vmfKJRh17PIXGPuzdhNofH80ymq5aMoY+AtSmjF9u43rRKaeNVgsy8MTLBShaO3an6Bs1Q
ALLR+1x8Thwh+0vesSCRTqZn1faKKK1Zx1lKuJtIPxx4rUbRKWxk1oYIjzvulKKm3xXAgqzuuAAr
zcNc67VJtWAbszoF8ZnzjjM3G3SssBiRwBXSPE3uqGoQ5sqBBZp1qti1vuRt/uUoaDjH0FoZHwLX
+/Zhw9fWb9JCBK3poECVTcqW3sfcFfBNnruQag==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aEdtgxfF5DqWViYScR5Bo99xKLUNQgRiZsz755OehHv9jTAW50sgdEWPVANfQF6BaZpfKzI+SCLZ
QwAnXibobMuez77/f2EGPrLonM/QKVZd+zKPSAcJ16EbDA97CVcYHuYkqc56s1Nm4gGkr4A4vtjD
Br/tif0O7K+IEHA0Q587JaVR/T6VCnbvWo7aaE1LW/tH5mj8vQiHzckWXTBaHKR5CorpnP+Jz9FE
w4gbA34/gsdm1ZXSEs32AboKZjjnD9VA79SL+2d1ZhV95+YzEvc6zb5EQ6oKT+BH1uU3fR1uTV3U
YGgT+s3RufEmyw7zyTKWT+vYe8of4LXdclV87A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lG8X6GS8OHba2k/dKrBnJ7/ya+XKpmuU8luVKMKBgUtp9/DOTd1pAOpxOsO8bq77vHuD8irMFRUF
Io6Z0+y+YyS7rFwPTEFARQPFu0+B9iRXBCeguTtpO5KVFD7MZPjMEd5xeFuj7z0WyBLsN2lTrSeg
BfZ9wT1KLMDxVvcAz+w=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WPmnyfXqCN5FkENLgZ+PrVqllbX3cIwFxLUeEJI/NyfHDl+Hr1H9hWl++/ppM8Mp+7mHeowH4Hia
lT0TS8kVIBBFSxxV+thgeKoQnsWh8cv5UO9vA2seLcVV2OwVVcrO8n33Zn9JgqRDXh8acFxXVnuQ
PGzEa40B1zXpQztCsiYp+ni4Iqs3ahcI2Cv97CU/zB0Z/ox5efXZjmB8r9BgVjNcS0T49M7cCe3Y
0l/bmxL5s3SexRYue9DJBy8UpLgNes2jFxYuB6eXqGX3sfqkmIXRoOJCw9Lr+MUsfEebY61lUooC
iEovEuONuN2btLKcNyWVKmiRneH/cj9IbH3MRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175280)
`protect data_block
Ckn2Q4cPtcIHMY19b3bzi7quaqOggS62C/x+r5nKw/LMwj6dW3VkCtSN4+TFmGEcUJhYgTDeEhQr
5DrJYtRpjWvJN0tf/QaM17B+P6mx+/aZEQCGGAholPApAFwofpX7VFIvFe4JzSJ5LgdEtnFSn1wL
gVCTmWMJFGWi+C0LHXnRYHhcHLni54gUDaCQRpvsViKqimDvQNDqin6n9YpP1xPS8/d7AhOX1dCX
lLAE8Ju4XbMUoyXPGbhRGWyNKyafTAqm82sQtm0FuaO1gxqslVXMgx2qGa9ypi4v9vn6ErBQjkeU
1xYAkHyrjVEi3S8hJkuEc47TmWOs/iPwUls4QAVxmtgN8RmVYe1ObDMU2Qw9oNHf8EvZwlcvRrTR
LcMrv1vVKgZuUtgYkfHHbuTDkZj1IYBi5UQF/A3i/ENUVBHFxea1EdQe6zk13YtraqNmMMXOemtJ
XmhML3Bji/Uolmvwp+jwnGJ3NlpBIHoIvhtyj+LXe/1DcrJ7T7FO/3oMvn55kmaFH1p82X26gbyp
Nzcuo/EBYdmFKRUQKP8TqDjfEx49CQFyt06SCyGRKIZ/oJrb8xykm3AhuArj77YXmJs1edBTTM0g
wh3KSVHfFYLRPzIvntsnf9L/MA/i5y+UPzk35g4NwOYt/IrAPc/WrOxIZdXmo8V8uSquirFrO46r
ccqvgX4QJ4glDAyWLuO1maFJ8eEJS7+oe0t4DJ8FZjtXZMYK+Az8mc5yyWDCpV/l10QF1Ha2wY9X
pnXzBk2XIXXv9dccNAiS5+IGC2H8m8CSpcOHHi7UuteU9rCjRux93f68I1Nz3knB9KeI4LOmIpDq
ccWypa2Zn8cjjG3PDadQFCWzXceMEQ+HnAc3NRlJ/OztyBq98hh5EY2rOO3r3FJCH4lTZNJsLd7R
HSmJ0u/7obW4WhAqlO8GJgrD30P9qLPmpkDkmI8WP8xdIIO0N4usx9mUh8LWPLjPRSMiLS5QhcVW
hVOYkgyGd6xHCRwjIzCxao8WSMIo3OaSG/j0NUcOmhUL2/7Ebt8RIo07LQ22nD7Tm+ZHPBElV1rY
XrpfHTeJ2qWB4jElo0Wkx2Y6ChYiuv3FmJNi9/4Yb+GueSCwWPgdFeyHF/EJSBNL+7VHyvouCAQk
J7Hd16BNaq2o5RuLqdxTsnOOfKqsOuPBAFTwTvsTPU1z7spFOCCn3naha0apU6Qd9+8n3iYGK0ap
OBdSdKMkgz5JbOggUNIiDeoM6GguPhzlxqwFQM40EVBXZSkT/mlx4zMmlPsZNgmct2ICX4+r13+l
PzNO4nKxfToCWIpc8K+zzlpaijyOFYxhVkYoQYsBQiCdgQj4m3wLSrQ/aAolfSNfyiYooa6qcZpW
ck7MJXWQBfBhukX6nks1KgISsGTJGE9rjcZbA5Ql2ta1yXcLMg9RVoFq7jL/3wtWySfIvVkUHVoT
i82XgK1DLB+XqK/n0QNM6xDXqPZAtHLk4VG9iApl9q1kCPdMUcSur1yjmmXCzGQMp5ZZu8yH3//+
qef+LpUWDP090QHfaWHc569sB5YVUg9gz5A7kmHZWs1lqUqkObg/seRp+AXA6rVcFJBxw+LERIW3
wt5q0+7QkiOi49HUK/UTxlCNndoT4SZ/zPWIv2D/mePEUszOcKTndPby3knyWFVaGNVfem5oy/fp
Q2ubifv29oIOd3Rz3Ao8igDeblIeDnq0R7bljDSidwCpKJ3t8N5+GT3k7EkSg8Tf44d/X3T+dPuz
K+vPKskH2F7IIvYcYGjKhYR6Tiypzd+2GhNEx6bjBgo7c1JpL96PPWLNjo2CtGiVQmIxNqqMo0Pp
I7mBRWKICijXJjRR3e1QPgqpBCJ+zHUWebZN0D6w8WHYfWDdkDz9kjRMzTljYTm1o3VCtlDH5t9A
ijPIHjf+tasRSFKu9YHMp+F5pf9abWadCoI9QSvxggfHe/Ja1GNkxXxnaP+3CzMqARz3HJytcXoF
fcIGh+620mWtPj4L/b5BxDQxWt1bPDdjSGVLo1IXTSOcWucngFpRefreFMELTOR4/EWp9QL8udyw
dMv/S4+85bFP7cReMtIvX50CTDLTtRWzpbW/fsy0WpmqXf77xaHl9UR3IG2XqI6jETlMrkk+m6nm
LYxoxcjoKSmn8Smpfe69fnWm033QMgWZnon22eHJIYd5o+I7MIX2p6sQfAvv/N95GG8DIDv2rNdo
1GT9auhtM37AnikEN36umwBYn4FkoKHokvxx0r63Py/szXOSgBhSoo6fSBmiejpVPDPCajLQNwZT
gEbqrH9LXEbelGMg8WzTEARcxuXwpAFE+ld83yH6i3Hx3NU4BdPb+Fb4GfUYOGll4YpoyvxsO2C9
Ipbq12xThLLnm9nqQ4WLPYDiKKF/r32Lhjl6XwJ3fgtKOSL4GtzjQq5gfD0A1UgNcixU617Vm4Tw
1VJgWser+d/voRTiZG8xdt30DNAs/sqWRqyfKrKs48pq0eqV0irmdOUdlzH29DZQi7Us15ADfbkB
PuzI4EmVZuI0cI4h827fJyGn0oAY5aTxHwrh4QBJ+PZxIbjFcVUqJgVFgm1Hwx/FJ/nv8QOPVYpN
TzVITHQJG05x2JKKw/C2OyeB+BBhiPEwaNt4I+xrdHOacRT6O5pCx4lUjskHIMHsJ+vOuS3EBF62
UrxOM2JMCVjrdBIkKyGCldVvcBxxB2RondsFjWgteuspuua+DIz2BVsUEeQTGyGd1yGdzwHgRdAi
aj0JqeINBQSll+Mlh3Ul2YhzKhs9TeYOvG1U38bYH0zK/ymW71gqU8G4DwKZWxS1qOHOYJwjxuGZ
+tm+MDMrc83+8VFeE8fkkkFHK4swNY2dq5I8XIMyDDhfxOH131FFSDHFvZLjRB9VhuZHrXw55H5c
RR6q/jX2dfhN20i2MEGLI0qKyxFpznAt/b6Ljq+RVWpnvqTHwvs66LNVUMh94uZk6VFmiL4LU5PT
HZBRJEkke4T3DQhuitwe50zYcv09Gqy27SHSVC+m73uTynad1VCk57ZK16xi9M3Y2pntlsGZYHsG
hghnRCGcWNxOz3SZTuD4o2FauCydNKVnDwlVEctdDUy/eDPBXkIQONoaL68a75f7B2sRFE8mk+wp
lrJ1reAcJczUg7oWiuLAjYfy6OqOaGcLwah28ZMMG+xBzFC2J6tZ62nw+XGTfaJlurnKc/GwHf2J
TKHTx8j8HhOhnPNGWWkwshAuCTsxKXIEzFvGGe0tpg0ysRnMeR9kBdD6WW7uMRKzcjtuAI6HAt0x
M39Wnu0fMx13XBYmfs/Fuyu7ytdE739prOjqqh+xRdIV0RBXLstZtvhzr6ljS0rinjvaPE9hxSru
pbqouGx5h0C9iv2259G+pq/NWi9Pa9VSiP4pA7jAtMgyoqmQ4k31IY48u+rjmsd6ZWe0nByzDOFk
4ROupltxhn3Ki7zG2mZWSO2fLuVD2iK/LKcNLEfiPRdskQY653LjpjQ6B+uBNMlGnS+JkwoFWbf2
xxrvflmVoXaMwRWTp+L6E0Edtxkw2gr8Q3d0DB3P8+rU3i0ygl35zTXXrYa2NJAkPxVjJJnyIYoG
ARvoxIp8Cn8BEZZO1dRAUug+ijb3h3q1ZlFwBTyC1subiyoQw7w55ucRiFlUgRrgGUI9U4szDaB9
HBCyJrYOiNErNR/Ly8Vm3nHF+dhMML2hf0dTFHS7H13PBusnsoOhD+atPWoGuZh23VLZNFUa7QB4
kWTTT8oEBxnL7tIkvDn02GDVkUnKWKGlZ6teXhGf+lf7c+OTg+gIgjPCo815rTs7iptdo40no1TG
a7YVSr/LwpZw5lnVLX03s0s6NIXShJUwfeiUZcsD94CY2AvsUX0rv2FHyiQzecpeHvULa8aWzQpt
hB2NQZKDYTR46XFi9ayxsKoeAjODc0GgVj7EU1Z07jWH01imk0awl5m9UBj4iPWjd1tOZUi8rcQA
x2pBq+HIK8ztfNfiritCZv92MIyY3V0MQXYh/Qh33D0yzXApXBTgyM2d/vXEKu6zl706HjZgwV4p
mea1cHNp9zoMYmrn6YL7OVoWClh9WQmvAtO0Jcp4XyXetzyFXeNTNqh9wcjV+5UKYeiuSm2kcyQN
sQ+tTJ73pdxltQh+2vHbOV9uGqmDbwHzskEPdGmx5eVmmnfGGfKMoPNtAbRW6jSUDm9mH1CAhvih
voX3e82kDTXx+vIWIuGdM+4THR9o3+Z2CubphE5t7YuIPCQzwibf7GgfHwMxop6+qkLoNryFAVhU
2uV1cA3XWOVCcSmS5V41PoSd13nmZY+iv9x+/GESxo3JW2LJreMs39le8zAXKkAq3q4bdMkN+Ewr
tj/NnasMg7h9dJMDN0g5BKAXG1XnuftTVpfpN5rYOKEiTdziFHqCkdW4ilUoJhSShozuQGXFxhax
BXScGUljSgz7zVI3GHFlk56OUAJ4B38KTUUyhxpUefQNj+fSb8aGvX9P8GmyB7mVm8AEn6kkcIXG
ZnBi5WRbBwko8lXG0rVHJLLz/f8qv18YK/WWiptzyPrC8KAstBoAk1bpSvbT3kcnFPJpbdtCsZVx
fwTh8z2OsKUiIds0nGOd4yndhA/zZwF1dvYa1wCct6h48T2cRW0h4BtY+UFWbDqyyhOZBTFbfKGX
HRWwPKXrOHJk0hKpolDy4zOOwGNHfwkJTVV5vIPIo6JOPlev4rHY6RYG9k1643AL184L/PtyOXIW
c8rH+iX29G6/poKwBWPTP69h+bD618EkEMBkRMgoZBM50jmquMQv4ZEib1Yc0xK4f3gXqNTi88X4
pPs/MJjrnRrXBEygtJYULxKEiIKHvXf0F53BGyv3rVQoljLhTp2rZBhaV/b2DgZcTJtxka45Gq9L
AhhRuyioTtEUWofpYIKFkIkLRcqDJPKts92AwjN84Gi53ALnHrvPYdx+xyTHMhkHTXIDQpLYDMI9
9oxtbrehsFodIShP1Vmpzgo27tlWUM2kf7FNZbnrPmMiEAEcRRbqNK1BPzk3YoEK4Z+WOBV2DVuG
ZAbnCz22AcpOtgOm4piWMeVb0v7USQ6LRrZ0SOjThyEi/OC9t5Dgh8iIClinvIKo5bSHnhEFYNuO
2KYYTU0SPfvbF5wcawjtDIZgFTM16v//404vhBrWw5gOcODwXpO92PhWYRF8mwxdfvmgFIq0lwEs
Vvy7Vq265qJWbrje/2lzCR3jvmZ6QLS/nDezvEjoJtXNfJEFblcSn0hc++DVJzrNmt/GX+kgQ8pZ
AlKnqC6/jK2hXrhrvYK8gbRoi8WCoIdLNyvl08r0rXw0b3ZZoDSWOa+0hMEW1lvon2My3qlNwviX
J9uncyzHa04MSGr5C4BI/YZT6FcCLbjrfmRbMn2LZkbItegt3iWbcFGCCMoMkLdPiZWDZz9tuQVK
lNBoySHJBm4wnsD1kqux/h4BCywcsIFNGyqxQWUIeU/ltlAKQDcDUvNsA2HMWgejDec9YS8+iErg
Q05JbzMPVdteNclIbFB5uGbGiEDYnZ89UKwzKae4uEBFAkbrgccyNA9kQeA7J87kmdIws4ICQVNE
k4hoMSjGJ3FG5DMa+pBkUMaChHjCiGsCvTDQC9CdRuU7er44b1VUP0mfJsbEjqCVSXw4ekmI46DN
fr1TijJH/gBNKk2RsZo/GDkmx+aW82AwnTdbZOXSjbl/dpRpPkjOV2Zkcl+uSS4PaEiagcXAhbAx
Mn7FCwAOrL3L3R4UwdpOgbvDWvZ4cHV67IxD+kgXVL7G9ggHMNSuXBxi1PB41oMIgOW0Ok/n3lRE
jViov9PMQBC2vz0ydK6WGI0Je5nkIfLdbwHjKtjflDwMnrpSmaQ2cs02THJsOVxkMcN1fBVQQ7Gw
QLprgP+VgJ5FnvV4wl86/fdaBFf8w7yyyCL2oQ4e2k/b1pchzZJwU2PVGiU/yFC5RQuhpXPrUV7e
3AoUlgAZg/DkWpvAxTfBPM6F6+Zt+OnpXY9LFe6lSIw6PZF9pNsmhuBmuxfwkhmwjAU7Fd90XHzg
mKK704SYZj6JPLOfZELFmN7W1LXQMJKvAY7Jgs3fOSpVL2nTdk9t2SeGatrSeVE+RcQcKz0+a2Aw
YxNmKyXSwxVYWutrXgcpbdyT99vJgj4iGunxaItO5j3NmYbGzOVwixJFiXdfY/+un+VNOCixettk
aMCwnm4jiiD3x0A+hXUNQNFejfT8Qg1MNK1ZkOxxqC9h9k5x4ez+Pr8BbGvO5e+i3+KGiI5soUPe
gHk/ulL9dDYt4CBlkZPv3A6aUxhgb36+ADc2u8op2+thAtnDu132VNRC6nShkkvLNuTNrZRE8nkX
aiT4iMilIBT9GDI+4JYv+2NT6zndkxc3hEwYSEc/YjoKXyjVMwsZII8Ra5+UbhgWYsvaFz3cA1k/
lyAQOCfBFOClh79XInPX3wcY9xx3+7lHnwbTSyQ7nhAc9A1RvLs5pNH7uyk15KwsRa2e1XsO2KmJ
e8etP2WjUPyztO9tGZjtYi1W6Ny8QU/IcdNhtk12bcitz8we7WMljOttppJyRxSTG9Apn7ND+uJ3
YlJNvHRHfk/a19mNVM6ksGnuS8qGYchkQtQLyxq0HYmfw55kA8Y99MqvgOiKCzlHXLq2FQwvQ3A5
rkKW+xa8/Lpbw/69t6ZCJlrsMSTt7+2aEReahGOwFdoeeIxvo89803cGnBgDPdzDlVp119JXrx+6
4iUm3vu2HgmzLGukCvX+82pFvjZ7NSUFs+RXrBs4RhctOUzGsU/k6mvx77+1DyJJaZAXb+zg2yS7
0obvq6zSpCjFZGybzfF61D35CUYPWzNEPujzorr3HskoCB4fS7FJ0vovviNchir+wg6YlPVzcHBf
yKEc+lMOmz4+dIcSWE7udm2UE4wnXbpDaX67UdM/CAnou4I48sPg2qHlxD0YcS+toIavaKdPzVIl
A6Xb3dox4CEbXOGRLVsef6esjQxjWf560s8Pah9ydXp89dBbMSLyuPn6Y3s0BhRFQlw1Rw6bD1fm
vej1n/vWp/clLXU68dJDTtI3FvHbq+HQp4HMs69X87ubRQlJcSXa0Nt5TCF5xGKk89gj+U86pMLn
xzn4ZMZ8YGh1K+rwmczUVuFcUt+r1WEt3Nrm5Om5EGm5mSuboWQfQesubVkE5qkaqabzCixjGCom
bmfhyhp/jaFibTW5odgDVPhJUmjYQu6DZfFUnP8IaYztJMpKIUJeOrxF6HfyKytoao6BxqTaXWCn
UswltS1Drn9EKqeEeGNkVDgVtZa/jP0896BvRasBhuajhkS+UeWxsjmWCZImvOe35zi5JG9O3ltj
oqxrtwpB/ACkSAms9RZGS6luUmPDFglhg4J4Lk7OJaq5neb8nLsfjscyjQeNkWnBOj6gKeekMVgJ
/m2dZzuJxmkSldwYAq7JZ0pQV7k4CtGqc22srliPsyA3K4uofgBDsIHOt7O4MnpG7rruRfScijEN
6JBaWd3lQJmaUDb1oH4PFRdzZ62r9LMpzuRS23tCLQUE+JW8Hws79tadEQ37hcFxvhYQ+PaMCFEJ
8581+ZOWriN8RRU9qBHvbhiv+BqwjZ27BP6SCY/0LQfSpO6nBMhaJBgtmT+mA4ktzQ4nZs05qySw
V7dwonKHcb4FwadDduXTrY/r0iRzRlGXcqMbcSEpLhWm457BOcP5loDdAqR3tNdKhtC3KF49PaHb
q4/yWWBovSL4zKFuAZm3JRHW0SBuGGcuZoEfsHWUWbr4isKB3J24mroJurki4zI5Vrfrh10QyMk5
uSkYajGzTPGNcqUz2sWH3moYfCQ1PWMPgIMlPwcsY/M4ESZ/EmrRI5T8RW/MShYelOjbf60g8Ck4
9iDFucTG6ZPA//24vJSqi+rBDCONYYIVUBFf7qlov4l9iB8kx0pyLtffGN2p3c4lMQSARfU5qN+3
Y6PwYloszPK62zv+50jN3wUrBp1dhHJsBVYyQUyHV67FPkY/bRW716/SDxaFesRHIFfZ9U75OVHp
sWnBEWhdAg6ydHa9aA7j58qw7mJHlR330+gQsTH9V+/hOtx/9+yzlISe+azddb4LLVhA7p0JkHgQ
ml6Ivxx2yp4XvKrVMebsgw9nXm2sSDmv+9k2QuqOU2UOLCicGXXnpfk8YH/+8RHzNLdsKclKoUYE
SCliaj07wMGembWd1iDNTXFUnmI+VZImTGEkS0XPrb/y459wp0WIT/zQdpNv3N6qDreagDvxiJE7
t7bJjLh/ZCPB6BWhQQIUHXnRWm9g6bJfLQJ4qLxODIV4kAXXYXr5s+UTP8W+oNhyS1crlVSbnV4G
xkZ9In27oo+aXdTwrPlHMYOyrc0AKJ9f9z9Ff4sHYIjwcyfbVvvdCUS1k4BXj+JINbVWRHJN2+zV
zqkAB+jp8clLqP6FdITIMGwP3rDs3JS+Clzr0mdp+BwE2l4hSK0yQ0jbAEeUTWg0VRKBw1uxcByF
Ai7sLqqx0ToVZlr/boarPN5qzB2VRXazSBstnRLOvxQTkYGazy3Py3uw1c3n4lCe7XsrGl6Vq6QX
0qLa/oCsUX4nUyBgASrN4cEOjpv0qGLnDYfsYsKNVqkn2yHP/G7iiRPplnkHS/1Zi/TzBtZLwZbV
ZI/YArcqabKM3lYY+C6MZUp0y0iVRydA5DZiRMUOf793u9uUzJ0nX0XkvhswvOlpBJKEEGBv/lLS
X+wqhCNCVVrJfo0ml2n2f4ZjRN8nxzjWSJ7I1r2mJq/0dR8+VzxG+1iIncoLvvf31o6b5ETSukYP
f3Sc6hRzAaoUq6fFkNJLb8OZKX64BR+/Baz4Jc2vdTKB7ztMm1gg+Iq15GNjDJrsGK4r1YFHzRsX
mS79LIodtq2tJ/+APR2JUJlFIkrerwacRxnjsUL7xJrWiFk3q8e4VDCsFL9+bHvALLNP3yGEL22V
dbN6bqVEpoaKQwj7YKAh9xL41QBhrhepg41JFtuW1wcBqACM0pljpK2KagBluw3VKnfwSMj6WE2i
Qy9daWBVbH+qJx9R+P0AtUx5uV/jZ/OrJi9/A5YExyQ9ty8kqCeNpLPHM1QKLipiIUfGT8YItHgU
b0kimkxM3WAjkAaLAYRjuXVzvCfAETzDGbzkOpVAPRcCbxqSwsqoOTEj/TljB2jq58udUO5S+QNK
LkwZs3b4IqyHhi6kvXRHq6NvsU1t2kbMbVakLSHot5/EPUMVkfnvZTA8JNIAq0SrNtEMpH+TL6FR
WpHS9gYhFQJTekbdqH37TX2mNDNC9dw/8WJaeul9oXB6aIhftZPUT4c5R6wRv+AAxe/OT+tt99Dx
yt+LMXBXMjL9kJkLIoRzfs27yRPbPIwUcXOmIUX+0IRtPjagGTSFKCT17Nxoq6nHFYFNfXaA6Mmz
8kThg1z1LLYRxlL/gmLW9zFQ55HipTbLgyGploBnDoaBaBgOVsmaDQZFje7GXRxQnaXBsG8GbGLR
IQVVtL7vvP/MMAARiWOZoVaWewTtGQ9DdFhmJmhuA4SV+xsKlmmbZlo3H8+SLC2I93Osmj70ikAk
HDOoSSL8ZhvfAu2vChPTP5mYOihK+FbxnePHA+JVW4+bJZoauRL0/1SNV//FpBhAFrqfeDbKNker
ICyLzQ/oz8hF8Zu4GpQvlJgf3mBn58MZdAufww33Zo+S8aoKqP29j3gVGh4XvdjP0uKHsRXv3C+H
D3clJWM+4ps4ymAkjWfe/ZkSnPgHJoLNqjQ9nTTZb/zikBtg0w8+Y0rN+4f97fYFifwQhhOTPbYt
bfNGPCkH7gR3PkAtcvTf5n2DlnZBg81eGc4FWlOGliA0tzZjoCwL/JkvWOoQoQyH8tWIooL6ZpNU
lSI62n3E5kzMy25G7a0QkL1m4Rjvx37aiA1mL1miTM5WQD2Se+e4UzelLuU/N5JTrwqYM+08m8Aa
zetDIR1u6835BktbEDSgcC76vYUx6SX4My54jh0qVYyj2CKlarPhSJwWyK/jhtopSs/4syXL8H92
WodtbmD51iz8kKTUIa9qFxp96gwXvOCPGRoe0eaDz39Ot3xEtKwEuv1J/s9d+IhgUe0gvvS6SJt6
d0yEhjeYK+thZ1VnZ7LNmRYKwwuyUpE/FO/OqY+1j/G0MQPuDrGhwoEopIr3N0xdt/xccuw2Oq0V
xHtPKCKJCjGqiyrzLQMtDupxNX+glrDz9alysFD6u4IzlAc9RFRTmHj3FIFlq2iWvFNi6zysilO0
3FzoorRgYaA5tU4KVBsV6xHi8zraI90iwlcbf3CeJyP0tqvXbwwvFyQT/ViNsDfUZGjwjk0xAsYb
7qFqKYKFPuTlSpi+Lm8U2WnlJP49ZCVdJJC4Faa0Pd5m5llalkrqcpm0ekWD7pYTTTw5qPMWMArT
Vef4fIMVidMHQe9laIptmMs4TZsbbLiPCNSbmzgemXOOsN9Lt3N1V7bYNN3DpNQp0MdBxsZjYggG
vcarr9TYZR+sKuyZtC5nRMnjcwV0I4Ib8hwUGX355g50G5ndrlr9izVtuQ7DMRCmbMgGdGUF8cAw
HHBB/1iNgtkBfe4jhoh+dWRf41G/Va5vsKPJjcWNVTRU8o3rBHO7q+2Qq49tbcrFJVgxemgbP637
c3bJhMwuEwkg6z+FW63y/8LNN1C5X85GXNXnb6kQx7pjxxAu2tsWg0c9duZdk6pJJ6jAFxlP+6MO
8N1EuSZpbjb0FIT3EYl7NAuTcDYNhi4PYJBjKUt/yoWI9D2tBb4ZGB11Xuim6XeefpX1pJ2yxfpk
cx7lS+u3wxcz0vUV5M4J1UTYqTgGRGmrxY9+vUU++RjEOTxl5r0OqXOTpwKecj6XNY+m+Z8o1CNm
a+PXV5NVRzJ+hEhewemZJtdPejhZeRtPMpIW4sqI/E+AGT8Qhl5CWkj3QxfSA8G8xEtXSd2/kGPS
nfkYVxF9hknOSnrcWFh4XqtwZWYGev+mxWFWiZwWCcSxnhx16ZXdI4lXbUt74PJRC8s95BigoPlL
GUt8B7shiYRPkZHLZlxpD6BuZJ1o+iv4S3AReNyCRt9vTZ5XzY05ucsySD8rRNBOBbyDRd1w83w9
OUPP7YzdJmJ+RlTfgsHoXRto2J+DjnGPKxWqVNJeUC6msO3vE0GYS0dHZPaxijFVsGyvc+T9Y62i
D1MdBsaYTzxv/SCh1Ofn7ChW6z99PZxYmIjCqP8BAZkBNNFqifflGoWSxEuKBQwnSAQDHWuDbESC
V+w7NhQHXlnrrvdWcfJQ7u/rZxe928c6rjTPMBol0uIxYsBMXH4S5ggfNSRhFHBX428Rp2dWIq/x
/VaZUnOEzftomxYCkL3u6WCODOs9v41svFl+PbDE1fq85/LZ5mkvkWtbftXxxD466+2F7MOROZlq
v6RIXkYvR4UW0z3qzEb0tokUQreNNI4S8EZ32Y3K3zvSqpd1SbtMd8prT8v0PuUj6y2R0Qq5wRmK
KDWr4a6jMhaDbuP7WZkXGm3ZanVNP3Lv3oGEPKaItUBx2OlA2m/qRbG+Njd1QjY+Nflh4GxhzDE1
utkwirqzcD5LQ4GSyLjnjFBxCpyqVsQrJV6oOfdpQXxeMfoi6XFLfMuh4vgstinpRl0EVtyNns2U
CDW7fDlimBydvpTFQINT0TZZpXz1HrdP3GoUreNWTJ2G4H4WVijOeb2J36OaW0+hm8CKBl8VdJAR
aEcioay6t8pkMbBcX+629Yq7eUmqMocE0bm3OUVkWwTeUK1h4X15MaCuSoQfaPIKSt/UmxltdYuP
8USQamN2Mff50+0PWtxbA6Apetn5HD9Ji+VY3zpOLjlRFSA0qQeX5DQaPc/UbsjUhDQGCavbOqIw
KgymGlwiD7PsN39p8hno4j9CyXDJXhay0sKsWKgRYiChzV2PIhhD2MOZYdXliB2qEKvtWbdK48Wx
RtzZ4QhDKXk77CL41uROVHXdY5mMx2fYro3C3j7qImjNI89xdtNtVHYyyx+s8B5W0U98ua9OuWEu
Iiwcfj4G0rmeAOe4ev3kMhkPo0xffKXEVbe8fOdselbdIBplXjfaJAdh2kwU4Zl0kaT+YPJ+AIJZ
hZJKSK/HLnU6aqwqcsEbPJN7MQ97a0N2zgKnK+l/tsNKUoUIMPMhbt6q9qGj9pGHcAqk5tM+Lb/E
8LmwgSt350xPGM7qOnpxut+AAieoI8JzAQtl5tYo+PL2VAzAlzmzP/HLqsyZPvN/VUgVH0Gtk1Xd
wRxeGJzrhw0H/fU1ttbzyRRUNxhXxsGgbzkbqHTXR7uub1xJNpbmoAEJ3oD66sFBt2OYk2DPTnyd
v7LAQQZ33kgdox1zEr1XrSzu2OCwZee3naOtxdmUAwj5cGQVppzka5RkFuRgN2VglHgneaPM7H80
Hm2vIQeonQ6lggnftpyTSTyF4tdRCEGH0AoaoqhK8+1OkQTSxfF//7bV1E8fFf58lv71mdiHE9uF
ZUC1IFYfUTaTS6y3tr15gqEvkzQyirGNBOBrI6QI2lsqYykCEb8PBd2m9w3cPkDlov4F64O9vlXA
uxczEODnB0DOjTeLiasaX58QKoSjcmu5/BQYZIdoxlY4VROEmBqZoEueaCMX9aaYinYvA84iOZFK
FIwhZs2/jF+BM+CasqyPjGkirvhZtIkFczEiZ3JkOSrTkzyWqFzu1u3Nolo+fnLFuEICoVz3Y2dV
c4x2PdQdqg9FiyNxAGnvQ9EeCNYguloXwIBL1yLicifkQll/VYSSjXbMRyQCl5G7ZzmCyNBYqSXP
gW8fmK5rLvogEgpzTmhu5gXMOcnHJNUVddGzb2yVJcGtWb4CIK0DqFUCXIShXxRaNBa3sIteU7UQ
hfUvP4URfcQ1RgYarV5wRfoButOzcj4JEwIan/vWzmb+ESgM9WQPMH1Rafhr+rnbictHoxsJGTUD
+S+5YTlWHcQAV0Hn/39jtqjPoYrz/L0rvdhoQC4cHiXsP9R7LLteQ8zVIMxzSC1UdmyNMMpGkyhv
MNc6jUcqakftrcxXja2lY5KM5ZWZvmKxDw0tN764ypHSjZ3im7sUq1vaYClyZqTRxS8ZY8KSKI0J
HgouCEZdVOxPxvdHdavgL7ojZ4jCE1VETRt6DHHw8c3qw6rfqdMPKcLYK8MD5kGKy4RreEpifmEJ
kKVXiNGrkq904aOcMX5cbUCR72TjHlKIhXKQIg5CtpApHLRsf43g2zmUjyu/UlBiYCHiShabMIFT
Uq1ADY5Oo5VXotVOovPH2tyfBohkVSV4+py2mEJBALw5wjW+UKpSc61xvNcT7FDN4Yw7yYSQQNQd
1+VEh/MqMp/2+yK4JXnU5EVEnPDtDh/MFmb9VJKAHfwfvFolFc1AthqkkTnfH9707W5wvVm8RwiI
By0pTVyMj/oX+tES6bE+Kyclms9Okf9Dnhu3Z3evvGJJkJvVB9+9ZpoqcVMbCGZIYLvwxjS6qbtf
xwe3yuYaEOnhlDEWyY3WupZr5uQ+z8bc+tFQxSa5YhVkDzvwHC55axIhgoY6Uj5XmUw8nfnmTVX8
jDSbe5RbIFOGmi1+C8C4CagVGZYOz42PZpc7Uz4SyrZXtwJhtyge0CaU/1q6PaSYP+bNc44UlEjJ
4OQHdJViDTdV5TI5dDatazlddrHQhY0TtD/r4expnDoBTP/W/2ZpwSLa0kmAiJOLPPG0fyoTVtoM
lr/7qQr7rJGNDIr2G3e1x/37UUCCjthPx6PFm1TK/xCAt0rnq/xC6phsyp7bs//spij1wypeRy3f
x9Lc8+nEoSY3ja0z2KptNqauJEryH4P35/icaI26+wkANcJys0Qw9DUsxgoxFPfYW4CD25kYVdVW
7/Pa6OU5vxAYk1MGSw8BIuYnyigCevRGgeRmUapXMaC6qtDq6qERaE2G3Am4FuBuJoShs9SfIZP/
ku3OZobd6jTeDQ0lKro4eAqVURIwwvT+cNeKTJ4icp4WJwU0rGP5nErnNbwx6dBn7BdA8Wq/6WwR
+rhEN7j8gqlJQ4/Jhedph/ohUJZFrPWvmDTMZASnYFBKS1vWJfzKBqux2aDdpej7DEnKeEkH0/+l
7owMibz/p8mXjSahFm4gepJKfIdbCDhE9L9nKsOTCScmKmC4qPelzk5gakSfP7nJUZsbl0FYa7w9
V9qJeuTK6aZgbTRCcPW2wxuJ5V69VJmOUyISHWfRWKDTXmi87xk8XspVoZDXKdjuHTJccNkvOpkS
bqFrxqtAhD27HcVyYDfaKoLWuvvc3szgZMfh0It9L5WU2SA4OiWilFvREZE2A7ILqbl20gRnVtQ9
MlTRWFy8S8su4jFDSO97Jby2W7cHwiVmPhDlJ+MsmnM/FuSpTp7HnorXYFZJQ3qgff1BMmcYLFIc
cEwkeGVTX7shJbmW5sjro35tiezB9txMGKapNPzfFQtChGbsyxmvmX90IiDT5wwJZg4hHq45/38M
Z1D3MyvyKVsjAezRT7W4gzstONMy4Ns4AzvK3p2D94FcvxCizAtjDOM7Uf/itDxzYBZ7jAYeld28
EyFC+w3sJ/Z4nqIP4N4KYY7fxIjBfMAU7ciFN2h9ksVKXv1EDA5S06fsCqDkt5IiPgw0CvDQV1t+
CoVACQI7OqJGhfzwfhtrv+9XCvdkjTxHN/tPZVjqJpa42Uv78MrKp80LLZgEBBqREAPfdF3ZcUn4
RVq8JwEsRhK5uQWV4yfMppq6X0NAvS0a+CTMhWG/ufpbnDYHHZHiJz60DbmQoV1Z+vtc+W5KTPTD
vX6TvvTbLsDdpCbwSWZ7W6drJ5EJwr08hP5mxtmeVs78cB0VV5LZXXSje8bBFRLC8BYKBr5/H2Px
YvG2N+VfqzeE8Ip6nUSltc0/xwTIie7KXLMN1TYuMHfcORHFSQ4V4yaReVY2Rp9meg0r6yOLMU84
rOewSZwsmP1flOdYTGiDSj8CDM2CqT4htLAP7ty/WQAeIfqOmEyi1FjBrJlhth9EKMD0znZIHuxX
gTWT468pXEMuDVRLR78MORHuxKsh9F51tBQPHhSbAuX9tfkMdwm5KJckvi1UKQ1qk3FroEclzNws
45J/J5zJ/CZfvWbYvxBr87BuW3O9k0F8kK7bQIaKrwyZt/8REk6DVljG0xXBrYALNjeTIrbNWxp9
pseSHayCbqgnwksSPN1FVp8wTLoOizvuK55JLmgjeBZVHNcSapUTIRe/s0g3Geuu+OMsxQJiKa+S
SB6+V5ONXaVnmztI3aDr80K7QzwLHSADpohMtzzwWBJ9R6PKyIEgfhX5niFW4ej9LtuE4EJGewFZ
J1r6OXr0rGeeZxtb1qT7KiZe0RunxDXMj/dp5P0mk6FR1STahVAVBmMoopho6cflWCTX+IuK8l4K
W4ux25OtmNEZWa4mP2GPSRt7i4gxDZxZgO9krHf/WYsU/25YM2djXh8gYNb+6pxpAWNE3Kejm1Gj
bhKsTs0rdOn2jRFvZ5zFjt1au0182nqHZx+DvINjpZA0s4Q2ekkINnQquJEZpDBz5tDAwoU0NR+R
zr72G4vbjz2PtFLGqhEbpD5ga0LrnxUUWHXsdXWSHgFF4dS57bg7kNbHfQ3ZYuzHisGM+IkxrShU
wXdeu7W3iS9vFCl3v7346SOYRRl/y91qY7HFjUDwntbvhNECReyZS+MTcMA+p4i3nJUw71MAV6MB
SDkfQfJq8KX+/rYVrkMzOXJbgBwh2osstU6nY/xJIksdtFhtH4u0yXRf5wCsSMhL7tqe7Mj4IeDU
5AthpBVY15oBalHzu5Gdd77023g0vd/Cs5LGg8is4Vc+rM9hee5N1KdQocSrROgPJGeo7sMLWy78
Fr56dvqUdoebkRQIIAdgR1xsTfJtwy4e2yp4nxyGNZsHuV2tvka2TJcXF4FvLTx18zllMArkio4H
4iu74/HlmnDVmo+enfPJVoFEdyh9bif3ztaw4zzemZKXMYkM7Lkc7YXRbv+TJeImm6xnfSSNO5QC
OuYHkkHc4YoKRskTipTMkGZScTQboABVHbDA5KTAr/znmhqGKW8zi8Nmqi+s71WUQMezPFS6AiI8
mkGo8rM0PcpO+asgjM8k7Jq+mouYsUebp2iIhCZWesRAmvIWMs3gZ/P57CauaiTrjaGUbfOBbZGw
R5HGLFsY+SpJyx3JVwd12RoNKcdMtP74dgdOf20Yhk4FJlPARAw29XRqH6sZp9OnhZEeTnic838K
HPYc3plLSo+EwP49QhtCgomk3QllVpCTeyvN3PwmZYrL7ximjOSSZuAfBatyIBoJ9fWamEUG2+ew
8yq1s80bOuwGshJr2jSTX1wRXIwWJAKcW5yeai1Ds1a87kqvHMP76njznNaGmWh7GxHC+kIACE0Z
RSZopIWONmctkWPbuc2SLIE+4dvNP6iidfcvwqUU+nq4ggBU0E8NOly4PBp0ViUDjRX/cdPDZf8m
M5jau9ggmfsfBeCijN3ArrvfHQf3EfeByINeDQ16PWhpBFfpvKA1o7FmaYMpwh06RtgKgD8HT91P
4w27WXEbjlx+CEO/gVK9lLEGyPpK9K2Qonh6fMc3WeoXtTHg9zJC+CXo/os+zoa+Q3L3YANIOq80
vO0SsEZ4IQoaQuG/nZcs8IpDAVYXNEXTDeA79cFENbeeDgMN7rF/jrAeVkjErB178dxQaKihH1d0
T4TpyYp2tTf5eUG4N1rfA5ZyI7caivxI2/5AEC73qaY3zcyXLW+5HCEN0x679DMwLnTpdXv3YNzY
ie4xrPhX4BzJWc3EV13w2OGh0f1fN+OQxhAePar5lqpGXCOpOh0k+01xYbCTPKZpTDfO0gw0ZBey
4qFY9EWZHD5CPYuTV3VwCv/h8vcTrpamOPfjZ/8+QH4wF7TIixO9Z8rzuqKjEolc/0Lt+uyA3B1J
ieWupTF3R6QXHUIOr4Da5arxQ21OtQnmqomqayOx7hMx+CD2UQaQDLmwd/xI76B1bQouGO1O+CUg
S9AmPELa5pUr3SRbCu0n3dE51mc3LZZGPJ68DS9WY+ki6Pp8zmUq/Rik2zlmxUeucGTWHYupq/vA
1mdmMfJvkQXkmN1YoHX1Tudr8+a1+pRztWnIdT7Dznhz0AUOqbbaVHDSib2GX/NWTm2O8Hw8m/qw
6tr6IibZD3SZCW4AzdFJYSk2qnHfD+i9PlEoxY2BM+wIbo6g+bkHuEZrV2bB+Rwv24uojzOooS+c
nm/bQov+ry/6G3X9okZ7dnHzNjPxHPEp2PxrhXv0F0DSEzBsAoXI5Xykx5xlYv5IhoQNESiqpzC6
0rWx+MYbukvyq7SRu6ig2ngYqB+qqcnktD50fV6tInjXQrPKPoMtRss19AeuKzfIRNGhfr9CzLOp
54ZP2Gu1LeKBqJ1iZHXFEq03Q1MoBoRdJbEtGKc25pkT2Gd0wqAvjuoi9nSQLBZUVfrBLlayF8z5
zIgWQUs9RF7wBSL5zPnDklottJEKj8cQronldv5AdwTqe+1O++L3vJeFbomh549yNHBA9okTGY25
YHSU5z23xds6DY9UE4dwJGW2Br1eo/4ikFWViPEpN5LgckK7wGcl/Yz9EnF1kZLYbQhiYfWNvOq1
KtWxMgjk80+rrF6VlDEbi7wSj7Z1Dx5NxsoPixBLAWjvc3EpA7v+/EBkEBsz59QIq+Nh2WXA4n3e
Oo+O5UA8Tpy+8j23tmvsaxw9XSv6udXO9YIHrKTiiV4VbGOeYjsbmcIVYbZ4P3TpkgxaLmj2R7Ta
o6I8gVBEx07UAKYmS5/ssk3vD7gkoZiZo3lb2mRhJpQloVitYROj2VNqqr3zP71HAFLwimNx3ZRz
2V42SVqfjeTJhUYlgY5qX7bAce0dIOyD2J6y0QoLfSdpJkOGR+MaEuULZZh1QWAFZbspgYNyHXuJ
vGRdl6Gyurm6ZwjIdP8CloYF7NMKC8QEps4HeScXQ0jDo8jLujzpFb1UeU4ybAZrZU6xsvvoH90Z
e2GA6X5W7rdw1FDzyL54HjLJu95w8eim8KRUfrAoglXwStCiz/ElMyphmR0IJSe/Ao7BtS0HDtrF
zuvRqZSvUh4TWLYSU/k1vPqL6dN/k9jfu7DTwl5GOmhIWvVqiqWez+cpJee/Yms0LFVZljq5oeFh
tiR6ayeZSMKVq7dJ2naEDQU9gwIF9c45+Qnpaszc1f3bjtp77AM/W9kQaqWlpwW4eMJl39ka6d0J
5dm76YpjdnaUTakOpaxytE2aPiYgVwW9GSmvhhExVWrOzlip1E/5NF7ZmODKzCPvjIBt3uTDl/7F
nA+Zv+lt4KlUCdqKksV9YciStiKYivvBsyiPc00OUryfoH01rBY0zkgfj8Up+dS2NbxC4E+VOX5C
fIycpr2hvAF59yCL3eqJ/bWXwFfIq7HpLk1e/FfdaFvsh1F/7exTsuHu+IsUGWlWUkB66/PgzF8z
d7+Rffr9SYrQ474Iyy4MVJd23lzB5QhiGpZOF5PZkYdoKRQiHvyJT7sO8fqt8H8u/yS2jhbBZos/
Waqvo/B5qZKjXXHBVmTPht8wGnUS8NAX24yWvDspVwlFcB+pDVUWMzRMalkzq5AUYXJQw62b0ApI
mkSqWLSSZqIisdW7n5KT/snmFnYAHBSoCzPH95kyV8egGUYpU8vLJK1R/X4WgA6M32y+holbfl2K
iPm1HM9dPfQ1F2QcRqmKJFLWSj3xtgDi4lFHxgNtA0KsGhBRUSd6h9wPWH+N6V1lAL1ZY5Zp/W/8
9razLHgra2M+XTbAx2knLi0jAAlTNzvW86qHAAX2Ix6WZEPl+FIfNs1tryOo/GjAqwp280Q/y5cA
t6W7HLbQ7HA5tI2nxSVpV0x1T0ocTN7RXeFzax42/UZqoKnZKN3DgcKLp5N6+bU6ogAOg8waRUaa
BJLaOUePIYdyhC7A/GinB2N4P1Zb4Z/6pF5KrE4830j4ZnslnXriXzIzBWGcEYfxSUeAUO98kYH5
fO6Ms+OVoFl2XbRkL2zyEJnTrODcEyRPJyDK8vIR6F9Hr3md17BkIZ1FtvZzUMD6QalEV0jK1DiB
v0KRrDTerHmJPHfP0d1Sm1PRjrX+FjL3z/VvCEvWDlFSyf/3C0HG5hLZn0uCwVXIXG/CdEa/HQtr
eQcYwE2JyJ9kS/4THDUzz5LpgpN0RrPjROwmC/SgzK/+e2fP5X97Y0xOaDI0ZI/HU2bYrauFxTB+
amTO9ZttbGCp3YERBwSJSNORP+d/bMhYZ1xjgeu/5RQVSWAkW31RvBo5XqmKBKvYCbGQ6o7d83Jo
IArexkzaVDBfMzNpQk7X6Ohbs+DwYH3p/1/S64x2CkCz/9DoBHLxHt/rUorWIX8GEM+O5DaOF5Ar
PJBuJz/p2jrhyUHq9SInoZ6YelhwZf4a0zcs0NQnlwsadh/cWKiFQv5VNcqsbJ5lO0stMJOCi1Qy
XWjFES0nUcbCcHQSD2wr6WonD5x+11c3KAhBiypm7DhHmyg3ntIY31/UC8MD5hXTfX/YSjVcIpnT
Nh6A2T5ENXzCfDFTIiji5yKiX2zz83DhFtdrMlFODjPOkhWNOsifdNB1MqXOLOAIIDg5sPSCHf+H
4sbZ/pO0Np5a6mMR91BM7z+sDZ36E256NHWgUolIkrODIiZu42kZxEhlS/FCRkNueIgT/9NFuqz/
1OdQ/Qcl9jVP+336oji8RwbLii+c7U3LMRqtVkW3GyNS/+Vuy/HQ8ZEvanH6WLD4I4GBHmxDDash
vdAos3ukCNJ7LTevG/LVxxsdNlmZu1Yo59yxzs83k094itIE/0S2ccCeX3xKa8tqoyyfzv8kNN48
hGFqJ6pMtvdpTc0MIK2sNsE94EIX0cX6l/qnW34ufeKLDmbF/QjLoljp/Deez08o84S91+XAWZhy
RbPKFEg5aJs7uGhu4wSyhB0VxCu6C9fr6nsltyQ0s6YOhu1T5rVrlZ25C2rrZIUyYKGeRg+2wamF
Hs+/VIcaeMgn6wJlhl10B2fhmDv3D/FsmFtXoSj3/+v1Zl/UiWJP+p7Y3UNCBxFvxASg/Jl7SgCN
AhMOVpJL2ozght0YBTptYyTWho2tX5hm02rzxmuQHbM/SxY/rBPmv3NJRB2aBTHNtIP437XU7r5i
i1umnCd3xHh5AECtH6j3ptA335Bka0jjxw39RHaimVtfy2psxKEu39EUR6hPZTYEy6O6pY1784t3
RU8VzkcECLtONIzzdPfkXqZSLnhUO5Z5+VkU+vVbpfKVaoAQa+fkJ0BQy7kNraVdW6Z82uN6zfFe
2DvU7F7Om6nrww0z348JbjWNAsWsESoSJr9mcnLDuF6SlXCq4I/bFsL1DWxIbiwCGz2jPqBYI3up
udodY0Mqj9VjBma0PaepnRM7nSITgHlS55JCFbQrPKEe0Ur/3ZWNH+4ZVqmDTCmZHC5hrRjRk9BD
YFAaPL9FG638E9C+W/sw7ah6FB2lhxDHfwQJ4XinfRU+IzRg1S/p4A5DvQsdlKdLGVwAtYLI1DMG
8UNYuFo+uuEergKulhc5es92iBMvSQFgz13TeLgxjKZnuvxCMSLqtGMxPvJcsrH4pHsvXNQs3NZJ
K8CIJ8NcpGl8kg79gYVmOX/5lgAaSkGb+vy98O56dGcbVMTJAx7jRVDZsqmYuhB46nVwcFb05Q8T
iECTkJc48OKbZyv7DzDYjZIaj0IB4eqp1j15hW9PAfhXC02PSZQ3Wh04V6y+UA7hNTEZCSUWRNEU
BiAyCnQ+h/Qp/vEo5JHjmJRVAJwHLN6jAJaxSLMVzc8EBRXyxtrb+jBA0By/gB7tYJ/p82eHLt15
mCloS2nmzoz7OW2wk21TCnMFWneIj8Dyi6b4meemEfez4cLNwnGg6my/h5PwJKURxHWKFfXgki+4
q9+0gUWC6FguadZjpTptfibEBrKihX2JHkapFgrBNtl5jBZBQS459Wn09qg2lo/LMCVt9D3oU0lf
76fLzcyeVjJOP+QBwFFJxP4yxx74K8Y0HLB6Qb9ZRYldwVA+lfbfKMItGl5u3ueGX6GcMxYbqB/e
hH/LrZSQXQtkXFTOlGz/QCcbKOATw5fl3XioAjsODRgF9zAy/Xkg7A5SqTwIdGWzy2iS2XrBDelP
8VHMk0TWHzJcchMTwhReoQRRTDhLyJkYNJ7BcTt2IPQ7DnDLZD/sti2oxixQYq6j17YNw78XzsWJ
r6cve/p5AEj2JvTMAJh64rnf9+W//guFYAxCaYiJDnG5R1bUZAbtdrBwAahZU8EhaXvDqEfiDb5J
RfaxT8wIpGxmLR9Sf/oNLPkB0eGiPbgxRt0ctO4l1gQzTu4v0BrPd6VoAdhKlNTbJWsRuajgBAYX
mljSHUYFNxG0Vx7/b5F7zsR24OU2dzFUzA8t/VfHK7PXXi+LiPbmHMwWJ0KO0yT//H71imRJU4fb
9ToPyndky6M5GEsDicNmUSGtGvurXDGk5edjNP7dZ2tOMy/xk9YwugdJ3JBv26lc1DWGJEPlFZ+F
uJCzKpPnIJ6XXFDuWbOPEG75HeHuNOb6GU0lAzYgkv9Vvo1TcJXU7o/esd5SFFvi/KS6QILKHqUl
Z5CgJo23iLyly4IYAzebfHUeykpXf6SElHI275aneFeblY94YWW0idW3kP9wjegsTPC7Qbpn6gRD
O7M10jXjUzCZ6EUz2dwJQY9edYkTvBIrbxbKJTcik7LbyIwk68VI46kI7x3AbRN33CcnoV6GbaSg
GKbY5gnbSlTqcUAzyO1wGSu/22vQPKHLa2zX41iJvDKbEtrBwRW03zzCW927WaQZG5pC3jHzc0f+
VDDv3kTqvFhWj5vvLmtZwt6uyGmnU8GRFCwFXFui79+/oqe+H+XTRNOd5stzqiINQSKIklL2INL1
31ai3aimZaGWPnMzM7WzhC3uw5nH6n2O5U9EmP/SswgfYBXaOXc50Dw8ynxCFsAPYNHRxwb3Wsfu
mm/DrylzTgBMqK3kUi5ogFo4by+EspdTAgWLHu/dhCXQLAcGGdz5TBT0eTuqkFEJd2e3dcptgnm2
apkPDUkUNibCd2RG4agNdL9eVJ7APRk47ZTsiaK8Ry2Kg71cZy9rMCD/gDWl4DBcdzvADjvRvOl3
b92zL9bXdmfNf0pmWI9LtAU1GyDjMZf7GCqLSihs08Xg/M/a0SxGVVsu2r/neNBdDz6/Ut7/fMJz
KnxXjUM7jb4b+Kz+8BIdkLOAfbKodpWQPVzYv9GF/gOaPbnAjVGYJvqxAWR5u6oB67g5+uhLY1yH
KzAAfKRJK6vygVpLnZo/0KT3gMFn2Nkm8u2+E3twRVcQPzybgBQFlOx3tUsjy0J+77LjCsd6eONp
+baAavrtghhQ5UirqYR+qIkOlNbKq/1ij5UNrC2O2ft0mgcIu60vUldfLVxa2waXZNgZeRntY/XJ
V+fVyIO00ZkpIo782/19FWlLDFIloZ+NH+AyrCKoa9FcP9u4yRs+zSQ0qSLUvBRuBu44katlAJD1
hFfe0AnjAv1EtIb+UMUiGP3hXnIwX2DRDjNzYQ9uL/98Q3smgJXH0rbX6epeTmAQ73HEUt1u0Jmg
NouqGTyFdXGJBjx9RXXsFBTfGTw3OVu5cmzzNm3TBCWKCZld6Ao82d+1lyEjbSsLUTbblBbIijEf
CGfUOtifEy+wNPXLimNbfmB8B9IukPOurlXI0BICA+V01Joazg/FUBx0wT0B+HVNZmVs1r0cT/g9
kq5/Z9nEM+WVR8S2du6eFs08lLf1kGC6fKFDh195xCGlWFVeQc9lUBBfvB9fOh+rSVweU1p9y1mh
Qd4hMehMF6/ZPQlD1t/A6wBPVMAnfayyjTCONKip4xo3TDWH1l0kKPf0x/NGldVXIYXygHvOBoKg
blmryUki1dndSdv3Qkn/5FD7JIbejl6YLZMzlAxyNIpnvrmn7bdG9CnphGx24ySMlCtmtlK4mdtq
LyRteN9oK4BwdiVC0YX39T7Ac1jvG5IVpPE9kb5kTpEABOVDQCU3lymXhwQ3j+TLz4tkMXEaZNPq
rwD+Qc9aqd+Uj6Hpz3jr2PwSumuFgTOXqrQqT4iPBd/Ep9QB7z+UVjMf51hXoEvnuKmC3VTykDmA
G6SGTWzBb4GibEeTBE8PbsHLWrgMWuCh1KtSqBYy9f1YKdfDZoGivFQSwzjhQ5cpI77CjcnIANZG
rofi4murYS8e1C3FvWG6MzykaeW86A69S6IrSxKDLxXV/WR6kC7Kh36ITMK2BSk0bG4PsMoxDZz5
IQx900/zhhQ6U+hCtqH4TYgwKGYwtqXUTwNFPXBvDwZ9SNZav9vBKezuqc9q1TxuC8h1CXSPIOLH
MzEKzCwpbRtt44fLT4hdN/y2dAdH0FhenEMPC1yAdtlWRBMsqM7YMTvAL906SPiXQugUkdhTfpaR
TCl2mWjg5vzxOryj05ck20yhFGFUKpKmriWk3NOvRawCKPAFcUdiKMeLGnOOnTOipZv9pZawuVYd
D/zunDC3mHqPX+OvAQSIMdwyebAJ5OdR7n0nvfLvxhG9qU0HmqnEMIWrwz8cPdv9k/p0cj8ATGmg
vtzDd8T7zTmV/Ct2zyjKU3KtTqHzUTA4PU+T0aO99aCIGxA5k0xRbnPN3rseOLRKRssGbAj+5tS2
Mfwv2F4gjfSqrsGC7/LUrX9SimdXSNBANMaw5YgUiLKOVEtOhctIuKI8adqUQT+uW8hyyjuFJ/7Y
rTchiJDAfsXyBCIkHeTHsKtF99OWS0L0An7nhpwtc5tR9Pk/0mkE6l3rKPM2/DHR2bNGK0lIO7ZE
83aeuHvq5EK8XPCBKSA+uYxOFP2fwWrh2Z0VQ2mPATvzur5vdKS5pLIqzifyChNc20XfpqOBK9TG
boZsHyUjMmC6KHgvCvFFsDaCDICd+SVeylPHVe70sqbATzQyd2THH59gHgzWhieCmoMIH+9P54ct
/XgswNhoqal4U/xhl336cM1tx7gUKCnJhamiwLHvSmDNdBiLEERUtU1SLKtJaDsRj5CPc9ZZhbfB
AHeuSndCA/WuC6P3Kvqh3deAkpzPAo8hRJc0sWlIGJF5zPCGtMw4gBLVCX9lsFVvzkTmcunRd/KT
iq0Kn+42KBE+uidKOfp1yfd6+dQlwkZCVz7K+F0E7O+neHY4Oq2dkHT/Ko9qzL0NC8VF8xD90VWY
nIeOOFgxVh2UO3KWZYT68iul6o0fayOEEGOu9NQKAskkxGTKp9Rt/vRytI5a3wa8Blk1vCXcJyz3
1G+N1nns2DmgivWNdNQAipkfUwIu5ybkmg1plPJgI65mDby30FbSd333GV6Hru94+DZDZgHFmuLY
dGaO8AgVgFMOePBQfF4PD0bo/t7RErsmv/Du2fpfXyzBupp07g2YDAELyE4Kv8Cmo7ioGFUfHjZE
Ntg96y5osP1L8BC8XftNNUZfs1tSyqFKrgxaU2hrry3O111Nx3U/9nhEYA0+QkQRHJiBgP7WtAsX
BL0CQx96eWSGZPtcSjuK88Tcx0i0yFJUlSHi7hmnj0m1BkFOwrwLO/P374UJ4Wt250TeMARpmtJC
GyIqv1DQYDdjnq10vhzOqUS53gW68EWyRHcT8c0MafYiv7pWs2v1Yh7kBCFCeN023II1YGGaj3vb
WYRBHKApKJVxDecWN+l7m+DaRw6wKDkDEz4EEzgOeWqFs5fJAAncfNJVbvdQ+H6QEJzYdWYcKFXD
WvZcm8YTIP2XjpNqaZI9PjGDmU3wklDfZ8GQuXD8blM17CGouBmSorTBa9S169GbR4h8dQuV90n9
Ob4TJEU+8AJ6d6eLJbfqQGQAas8gk0+G9qHHt65WIupEfa+VFamXU0Fsj5KM/If1eLVQ0NZ97aUn
ALHKBNAARIhqUk1FXCLLcoC3+zvpvaCIfR1L8QSPqNIbU7FKyZOcBWNHMZ4RP6neLG8t5qK3vx82
UqxNtE9iWXYsrmXe+C4ZoIImkurcniKvfrn0bvyhow99dronTEXXKtk9sZNRVPfU/KY/bKjSQTAN
xYueeCsS5B6G/VP5N3jS1jP2hIrCTCRp5hzyM5w6aScyDIVQcJrJIQBJS+NlFQKI4yX7JIQZ7vlH
ea79dTitR7U31YO6/RtrQCNE3iity+uA4atEhlsOaEkCdh3eG9WokPC6i6Ef0hFKq4HWusqlURL5
ODBrA3lh2x4zG2nHRUShOg7+huG4M3ftDMM38jQZqX45aZYkme0jpvGE9OM/ZAVLsQ5kijWW6JZ9
5vwVgVjlkAVIAhsCM2bbbx99dO7XOAmcP6cJ5iML4RgsCOpLGfy0CwziW0BomXvGnoOrb9IDmtiA
22UZXJpFLSWBLV/AZDbET3UA7wHmH7l53S4yyul+ynQbDA1euN0EvGoL9kDattQ7TG1m0ya4Nxan
hpCeV7ZtmnTr3ucIYULull7R4CEK01F++gY1AQNvMBTLY0FvNXsqM+gJ+iSdboZB48dblVFdSSua
uSQbQYOLOWissKWRsio25IN5SNpNcw42QC0k9ADdnBaHsprqOcRf60/Cbe7Frm5aEVaYBHZd1hSV
XKvay7Vt8NKqQlFT+DllVHavCyJClArhMmp5tEfnCslwqG4akoN3zvCGGWeu82vIw8n9FT5FezzK
+6ZiVI9CJTZbQFPucwp67Ou4rFTQrbEELR0ADL46KCrHHPnNXwFIA0KsnuAAyUDKN+Pm9XgZweCg
lwl1osYk1V5A1gqEAMQpeICmCjMT1oUh+4hsj/B3qmPAmrB0zx1m1rasMHIfoc6m4w0r2dGgMaDV
FvtasKQIza+cUQCP2FID9ny5QeY3wz267EeeBNdAXY+VOv78hFK909VxeI8CinmmNkyw/YhJYpGD
I7Vr0sK6IEeWEpFtTVkS2ntQL0nUrGiX+J+Cq0cQlVTPS8KAOClt0VkAAoU/mWChELVP4RvLDC5j
uoHnCtKBEeBQLkfXkvd0tTQ1C5A/n1n3kiQRhlCGBKvPK19AtMpNoCRGsAvPM0R2HMYQM+oFQeSV
KywLL9oTT5obic5gHLHss75sZ1aX85TpVDgjuJm6Rah+Kbh6hQXorN2IUQprcU+7jwDUkyPXVlW2
kg9cGM3YfrQ6IuerJG/QSM+ghBhKxIAqlJiIwWXI6trezU5hqqNx/I9ejwsYtYFpXB3v7qBRGy/Z
eb6C2tpPIXB9cye78UknRXHGz4u0YZAGl9Qygna2US9rmZU9rbbMb93W+MIwLm1BwDx6MIhzL6oX
uYKD2OgCbccObHAZ27DI4VLKKItfz1qd2KbfXD+uHKH4YV3w5oTk0bogy/tTeNATnz6zHJWP7/3g
JZvGNeyAv4NI912VIAQU8h7he58Q+5Q4q6171cFwvTHKuNz7aOWjkvi/UfT1xH5QfJLV5pkafGYG
G8cm3/0gq8VRqcTj1pnob8M6zuOh5qMqioYHN4lbWJKywEoQpikME2wW73+/IEin38DxY7XBUpxq
wo7MLjajscHN15csDZtWEEgfzSH0ClsbZOZTuh4ha84sVwa/JnHv3t6ef8o3sm3N8CM48cUljF4z
fraFh/1onihwCVJQZslrA4qn+xZNCXCSFeCwS1uvVAd6VhBD/0igDNQ9zaU9YSgaikaGdOHog+zb
1KwxXFVNYyONrgR9Kcf3Dvr7xJY/wfxHEzGY56poMw9LEqjr0IEelt4FkIQWuCaC4JFFF8zN4oKG
ll97HImZ7UlGtSrED2ZAdnAcVzoZ9XlF7SFjfcGK2Gr/32T6hJUC+rDdN+eGFhftGYjd4ID0WFzn
CX0BhCFzMylcySx6yfjWGg5p5l7dvYytcLJ8G9EfmKQKicu2U7/pt7F5ZEtrLP0LCVj4BrLo3AhJ
Er/J4Cnwbrv7iwni1Vvq1Z6QY+lDEuWZF1rtlkCV//gBBQg0YGxQU6JclGgNn2+plCI1eKF7Dk7p
QtiZxdHFugrS/IfaCJ0LJWhrdV8qPfWA2MA2qcrkyv7k/TIn7ivORylBphWgDxiWTXDWS/LnUxEz
WSfT12omYOjx2jmwmVLxi/zbMU5StGQ4WTbLw8GllKu06QWswX6mFczyHb4i0lFYf4FjR+QvZvyW
zDS0Xc3TVYsa96Pw/N7ZtevtF+aEKhzV1caXrUlqF/OUu+NFJPtkN2eS99jms7BsWgAUoVM5ZGZ6
ntNB+E7N/qX8qCQgJf6BaLb3N9X9yfPXhDq+RBIblVa/jLVKKjVUR75Mwj9c/Z9z8cQDoIEJopjo
WIF4fatGS8rZpUKpSFZYFXu52ps5thPBH5OhrLWZRdkZXNgAELPdc8huPADl9/jcWPy4kzDKOVyW
b1uVyWvIfRZI4zMTSTefYrmsXCTooZhKANLTOHdheLyKhRqJsRMfQErZLJt1y3wJkowDtgrlJUft
TS2G4t/mPYTx6cBQpV5Qv3Pg7CAIZ0IgwYZNUqH8i/dipQxep6V6NFP5dTgEBzhJC8yiU0UT2YBa
NhW8/rsf+I3ZT+S11uubFTGGXb6tuJNidVDgenZsZ3EqaEdS7sYcXrl2Lk4sm6QY6I/0neBkMN91
NDZFhgnabrua7kGJpejVwIA0zwzAhm5AoXwFHxWjQBximB3RnS0wvtt0ROCFYrTy4Dv2TEu4mbsa
46QTA9OoKV2BayvZVw7PfTcbBSmTQa3OCBbVxjPFHF+pPzoeBEwfuuZ6WmwjSz4PYgf8X7nlDyy8
rve6DuqwIqtq1CBMzyrOTp5UWXikvsWa2H28dUmzQG+XRQ/EN+BVWivqJuVGTkH9JFMT9vSrS1el
FP0T/XuxCRiKgvLvHBBk8fzPh3iCCzRkcDNuNqttohpL+vj6m5xefuWQ8L0Joy7K6e7GIoKm5lBu
lbvsj3AiLYijhg1CKGG4ie6ZrDp/9Y1kq8AR0+jcx5YbIqXS4E2Sc7wiJ8LQAazFG260rjXCMIsg
5kNe/S2mvPjgcLCVEKR2yF6ZgLAiw1j7rrNe+yMA8JyLt/J/Bmwml4uuocKq+IE79QD7PuXkrIdT
LIIGd2UgcBMhR8gFhxanqjqzWN5+WUNvakK5inzhsO82RFmVEyn0N4MUdj/2nviPSvdUgYj3OajY
bOrANVBz/JpV6LmXBaqaxVszwPv7OaR1Gr/pMhp/f2INtQINw7pdMxmpcGRF+spLR2jRkTktzHG3
NGXwpY1V6UyUgiasuV2hmRwt75+v8askMtU8Wfi3VWq5eSdA0EFXZzuoviebh7MaZUfiKd0axXO8
LMMPqNPgIcZUwMYXHoEfWt3XPW/urh6ah+fDHq6KwhpzVJ4k3bHfnWFXuJLTtPsx55UhL1RdZqcr
IEIthO3lTH9f0Y2TYDFqVCARA8v8c/euUUv8QB89ZrRHla6f+TGHBNR+zM4A9rzNYyk8l6G6v99Y
6VEtw5VDkHSTAAiLBy+opsXkCubhneCGzokWmigTGpDHKA50LSdvlGgyHKDh4SeSyM4pI9RAoJYT
EqUnAgHCGSu+wtlvi7ycpxkfqeBz/ohnqDCNWB5zHUp2OQDKmSXUOdgvU5hLeyZj2l41nEdqmkwg
il6d/eQbS67QoMC/y78X1ZmqDB87Ptyc6Ikz4R/uPsHHr2xg6cP59UA7u5rTMe5TdAbgna0rOW3+
i/8Yx++qBZ55AoGjrErfR7nReysJ1Kqs8UC+dhxAfi1iegpwSNPtWwJWN/Z7hU88t/vxXaImfAg5
H01cd+ASJouqqaWkcnO64JtwCMfCohUg14+dpM0ABbYNOhgqoCj1jUccDH1N2/Vp0had1L/1OSRW
HXTRKO+Q/XaD1OEDnlWVLr25nms5XWHdmu7ngSqiZQq58EeP1BsM5SbbS5C+8y+p0yr+zzrOFlXj
txOkFkrtStYCyS6sfjqpIc/N/wgFeAWZfij9yErGVgRz7gWl7ntGRhmS9TztVp7KSSOVC+yuA4yy
1D32YqMyIXbcXuWNq3mK0oisCdIOyYbyiI1i4BVCNxiV2zayU26MPOrbB80C7cWMricgMTDKcSdq
QITH4VwtnJbM2Bn9wDiEHJE00wpyyOYiaFVw5ypGjXjJ1zCAdoGheDp3I/Rc5ZUpQDkguuzScK9l
gVp2YW5b5spPbVxNeUjdvtBMq+yVLYaM79OH/uwueK+khv/ejZfUzMams4sV0ICfXslGv3+u54iN
RSzkYUUdedv2JDesfYFlPx3dbG5N0znyN3Um8tSYyMUb5ydHON9TwMu3fQKsrsOlEFHXqoqTDs0f
XlHg794cDqfsD3vU+bEpmQx9Mi+2pmvTHyGP8VpIUNeIslbvR8U8QJuAnaCv/puf7LRrgyXTf9EX
AnPM9nrIijalXVLanF7Iavr46p7w1V5X4m88mJRBAd7GZxPktI05JZcdqP2Eqn/emMCpQSGYckxh
KoRM6BAjmuAKxS3dhNjOxr4RBjyodEWoRhYiratZ1luPCLU0jsWcRMMS7PjypHXIXhRneTDUMljs
3Pr6w3MlrBMBEbUKK4Xte6PYtEMaLID8F+5K2eImLJZXNqg7hbQNpLbR+qHzI38z+GsgqOCbM1Tk
aS7u06+ZFEKgd64ST6+eNOSvvEkDtQ1bv4zapkHEQfC33Po7ytsNsabqZWWIci+r/yaEjYR14Mjx
N0wfVmdMCE3zLYzRqCM9OflkgssFYxt5pbOimLTP15frC2loeAf9DTHRZQ/e+Yftav3g5hxt/CJc
9IFAlCQzF+6eQNNNdBXH/joZP4PUSTdyON9pqlXPnfSBMZUPQjetjOXTb01+NlPfyW+kLErQ6B8r
Kq7ReSU1ow2pQMinyxx/9MtY9OY2mKuprXToZv4gQ1VH3MqKOS97GWS1ndkAyWgs6/WONlwuYZfg
9eWRvvIU39aM30aIOaL0AYm1pivO9hGRQGaZPoGlEbypWw5fgt/CfyL8O21f/Zjp14qKyeFp55ZY
C1KerzVM7NvlecgDb+puK0SpXk5+FEqbXwGnFpzjXPAZvY6GVGGL9h+eJIxuaoXZDcLA7oU90XD8
nGm03E4qUbVMc/iIyeS7lZJ4Eeo4StVwxE+VdQfYx1YgNCz+FxePNCI6fhFmoQJLbRVRlaJp3kJG
2VQEQ8n3Yhe7CZ5okSdr4UyptTAdn/Tm6w8ilWcpzMLmDICpvJOXIWaRqzb7BY0dGj8pBh2c2EJk
Xyd3vO6CW7DHFNg8xKNL13mxEIyxNDjb6xU32bCSv86uZOwv9Tan0hsJNSJsYeNlVvmg+6gP4Kyr
Hv9OXZE83XQAPUr2mp75wG/irlPoLjsakFElR33S4iWe91zEY8lAML2M/VgE8pERe3MtDLsnLjzv
EdLoEaIbrjWeyO1jo3PigMabTKFtsMy9yB3wKANRrWs+H//dlBSGXb0C98cZG0pnRBR8OePiSz48
60tckp1eFC0scC1VeaMt/uPaFnfpaoMdtgeRR+uWiYBbEOhu7+6ctUxdmaNFhCJeZ4PhE+1DFTut
IzZYnuCsoC/csrWAhe4ZGmhys2a/HLRQm2+Sk8X0i8flW5Xc2CYpkcmn1Sn6PwkdF977VDdQqvai
Ussc8L1V7mLHfjcEiYH+JKZtoBIU+0teiSrnp+iZ0BHcn+uryl8QTuHrZlv242lnfCF2RV5GG7kJ
dcDWQU+Xvh1qCv3YpXazkZBLh6TXyqXJ37laEiaJPSHDK0Ysm/IRQ/iMlrmNYicuOTjDg+MHt1ii
1yw1JoqRpNDpG0f5QXwAhOTwqNoHa0aJIlOgnaBLD9RPCaSo26B/LXREJQEaPfEnqjBxEaDPdK8y
HR2Ni1tucT1n1shzk237cJVrapfz42hcNmNRMmC0frKhe14auQ1CPJwDCbmKxEv6U9F+ziobGg9l
4fu6xRGjP7ytdQMPNSHTKv9K+zmdDt7CSBNlNd21uvI9IMS3gijmB0PxSLmd5jR/VByuM0XunV2A
RvTKxcOHlY8KTuTxbPkOS9tFznye+6282lExUxyCBQVMRHdwkr6E6XIuhOLSufaE7MdObUNaH3Ei
f8i8EAQOwpkLtT7MPmBZbfdUKTu5JepG1eGGsUAWVCeUgVVZExNmS6VIUw6FQXc7iPh24OFZRBL5
uPZr2s8dwAi/t3JzPhh1R1E57/1SmzS2zgtivlny1oL68dzyp5gaf6ccPt0a4jGFF6wosM695Ppz
3ylhTx29NksSd7QXFKnek1aEmID5RjjrllKJOjkxELInygWpYTVBo+G2lvrvVw+JFd9m0NfA8Zrc
QZG5wv6TjO1FnieNBMkQBbZKVghEaS4T0e8LTH9/b8A6oCzcAylRVyB1HGm2ek8Gw+kZTfkZa1wA
Xuurv6OaqK5RymHRkQpGlormbnL/ZTOk+o3i9xAYcw1YjFU8hB9sulGo/xT0i0yoZ9RCM++h6LFU
p5RfBSpJO1KJHyIS0TEhDjZQjoHyJy4DAP3E7r9wEBKV9lN/xo3+j33pJpzttwOiAM7Cm3TDcchv
sLSgnqCcbaawVtQy72AZ1swBQYOoKhOgEkRXQXq2VRqfDVL+RbouQAWLu6xFamzUD2+CUTK1k/FV
UOy27HPtgxAI+jQibGm6o03MLRiLQTydFViCJELsFckEtDFyvJ/qfmk4M+jmNfGxSAUJsdSq9Xxy
D6uAcT6jgHNfwJ+zPrp4e1TvzmFjaiP4TUFxGh3h6u/iTcun5vnqGSLBDqIMPrfpNkUg2euftQDZ
Zt7LKByEgjvKKTiRsWCgwtUC68SyyAJ/VRctff+5vHuvko/K9RXsEfj/EwrFgEODtbN+b4pQx6XH
WSBXO1Bi/YNfvMwH2v66KfWdQ4tuDI3fyqz5TUyflymKusZ8r8N1rsx2dUVzb7LKuzTVUMrlG+ch
CbA0YKTHoDeq+LJvjwkeld+9aGus5NkcMyROGmv76+75yK+Na8J7X+s8XxSthuHfjIlNUeVOGGsl
VD8I8WUhxEWKaQlZzmZKpjfFr59hKyxT0qM7Q+4XuJqS2dfmZClI7PRv5RcBe5yjxFpMI9M5Al6a
SrkXdoB4TyuRXm5tsXhK6tAzb+pUvFOwa+YK4Go3y8ii5Doh8zMsZuJbyc+rkl3MGURR/77S1rcK
K4CF0j08wKg2Jafd2RHi3zsatpk/DWkQ/EjFYxT+gUaIt80miwKoiw4twp7NSVXvqyNpcW/Vbor/
P9d3AEvXeKAaVBaDuZYzNPkjuFj2kmQC+KQ1E+Leu3g42vVA3dlKjFB8xzP+ntRsSf/SPvN7LDCY
SQgEubupsc03MUI3VP6wBUxv84tdQKf2jTsDxHk8LdlhJYvKnO1wdezUItTGWertwSNFuMqhMs8v
oLN41ITH6rKz/fUJ/rNyL/KFhQlZ373ueuY1N7a0igl6SJG8M9h/uwBxZYv14i9we8DOHsJskEMD
b2L92XtqABd9WpNUVZtJlBOdB2kAUV0Q0JdUFpEmEHxrg6iHOFGREbuu1sdJZBEg9cHZskMWtYTy
9Rvlf+Rh2Tx6nyT2mrS7Ad/ahp5tCK033U8QfQTfpi2I/uBkoBUu/sWtaf1US9cIY2d7Jyju6Vdi
vCHXgWQ3Stf6d/IcmxLj6vZuIiz3r9dWhIxq1NOjUP/HO6WPjV//If4N9PTvfyWahb1FztBB53oV
fuGkwa+nFnURyX4E88x7DS3dvzjZlWXiSFl9nBPDHbzm2SewrA/eCB9X0sFJtw76qP0WdQYAAz/w
bGPauKTj53g3xANijm7lDLyX5fsdVV/EJo4RY6BG70sAU2JKjbfunX6oq67CDRnDPBCpSv0hqvYD
O+kKxksaTV+sryKr8p1XT+0I/ZN2OKQsZtcDBwMFBG3kCKmL/puov4lHI/UIoaV/izQqwxt05fu/
6AvI1jG1BGXjQh+rBJP/MhCo4408g42W4lH2ob0UBh72BVP+9v27q+cycs05rp2bSGoQD32eGbil
MPDUgkYlNcG7Q7VuRXC97nuj64j2iMIoDHbyXvHocLZmr3qYAch6Ikcfw23mhHlyH//ocp1kC9xC
Bs7NWtz/VM9a6VLwP+Ww+ScUN1FPhX1Yrj5Q1oAP2Z554X1D+GguZRL/FsuRJD+bwcFA+bcxJvA7
CdJF4V0PbmBpalDc3QBbZKAdwYNPy/CtYDN92zMBlgasOlKLs0gnfUOCZ0oxkYLArBzMIWUBKPqy
h50Kz+IOtLe4DtLgVtjwJUQywy21iQM/5KLF1D6r0HvWiW37v7bnD3AMDLaa9NQGjOl+CMOH78aU
mHUwpDjoCssB6jCBWiKWLmhdbvRZNj94+BONR1vOn9UOxrPcoWueBrdczp/LDhJB82jLLknVXue8
JQE557TDA41/ykphRiBS0ukGZYdiL6fGTjAP7yn/0Hw1LwzWsEz23PFFQSL5f1r168brYtxtwy2k
NH2EdPhkvfjbCqcHOLcawGKqQHdZwNq/fPpTG3cYzcoGaElKvhE4OXkEh8AuDUGOwMOoDHAlHO6y
3B9m/8w7rxeLMjnsJj+txfIySlh+t7kb4Tj7wTWZRbqH/GfDU/exNsaJQ1fOJ4lWHY9xEEQQ+QpA
26bl863i4VuBdzHFYqBoAQ6yKH8ZLWN9FJlIYz3d4fuexvgxEZav7iCHfdCUgUVtW0QyyK/bA8ce
zGCceHyjRwavvOdmA/GMFTsrH7/mmw/ncW1RxiKKbQBkCWPNaebXC0JcfhgLodzKbENg0nEaF6v3
b12VGFNiQSJ6VsdiUMaLJyoqLwPA292M7nOG/sutESh/SmOO4K1QzvNGV373PfURfxY8rr6w+U+c
PZI5yphsq1w7vmouVUSXV+Xfibudu/bss8J2ExE+E5UZ9awWHyyFG6n2Izszxia8EyQyTsl9LX2g
GXFT3wqDk2giXQSLneCPPEn3FuDBekW0uBpzebpZewRaRYJDukNWS+EdLqOqkEhTVcd70tEqzf6E
liqo12KYMiwZ1oZ+yTZCcR2G90A7OrKR+pXCDrSg/KivjVJPgEE/YU2gDOE+Bs1mMwweY3VoHikq
FMLjEWYQBKSYzED1kpaC3N/59jpEYcZ6tlLCfqm7qr21OIZEUfV6uEPv+VkGanaAmO5XRnQx2fSa
XKf/T+uTP2SaMG5tVNVfheJTKmPXUpRhbLj0HstoaiCjNZ6QOs6MsTuaUabpADpqa2C6eUFN+BCN
VaFSx/E0Opu+oVY101jvAt4P3On/SYW2+KvyXUwJ5LxWFDiC3QZ8L3B6Zy7DHQOafmScBz7IjKbS
Ip220tXugBcoosfuRLolx+srjhPqbtQKzW255NmnWzs4RIhkdQeFq4yA6ryXVNhEGeJVGtvi75eH
p35RhTxM4JB0I7y6jYgfvmZIGxJr8otoKy7xH/OWBFwjEm1eAzS1wiyICEEEJDLNDqgugk9yeHwA
BFEiCNqfFQ3SZyDIfZZpynFjqnLz0TG/I0ETeeRondQEzi4wyxBJWjSlgookVmERJdyjYXUUV88e
NxA2wqXpWfC5GoxgYVsQkNP+ACWW9BtFSBH7/4x3CCbmddB/cbE+7MOxQWelokDuPWicoKCFZdae
Uw37qG7X2Cq8LR0PgSMnnVaa8rt10TWLCRjdkTpCXWFbrBYrcVTxUV38SAQfUC87YZpnGNci+pPU
y8q4hSW9f6HkUeZSeNMOKIkW9ssc7XGgKpoio2U5Q+V8rbdlPyMDJ8zmZojJcJDR/mGQV1fiL5ds
+f4vki2yYHgGmSbYOvmtwrifSOisQd4AkONO8j1BRV3pyvbHdkN0DqCTZHLDU89CG5y3XfSt6yIx
UYed0l4+yBou4JTs4uXHwEJARAqpcLRcdxY/PEmvLaNny251mDxVVsWHwvDVhJDwwj+UejkVb8np
3HGAiyFwGYTU4IyfRAQPwNHVHUTiBh87Nq2y70xg2VJ7jZrYEfNVBEU9gjmU242T3/cK8luYrjDl
WtukS9YhuyV2Tw4Py8S8hRM3p5Y/J8h0x/+A6vQT3P5KQnY8xvL1T1vIxKQYgXdUZDOxUx4zU7ZU
XmqWdTCuV+gCJErsp9lHaqlJ9dyx4ZCF4i/9sgSjkNpWdOdxT8ogwdwzlQV5xGOcVKd7Js4QdIwg
qKbZGG8AfYhT4eyZGHQYQSJs/vKp/XIdYISEQk8lsfI3WPKmVDG0smQr7WXwFdWy6Ma92qlf6vpI
h8eZ7F6VHwWneOc/5mPYmN7zdqgdhmuFxx5q9upA4HkNSmR56GKn7SIVPGTS6oblae499D+PWGj8
97ZOjiGZQDmsU28yqZMFMQfA5SzBiW6EpfRG68yB3jed7M47f7+bVCMjFMdAz0nRvy3Zi1z1+L/J
qn76SeCIiAAnzqKkqlG8+sC5DJ7dAXWR8sTyIIHZ+ik46NDAl5D1xB5RhVs65s+nV6eq7zYfJm7x
k5dS7BCwNAvhksDFJl9xFkMSFjraWuM4oJvIitJXLnfZYxU20FNJPlm3fRimYFzV5m6WePA3y6xm
Pe2+arxqV9fstMEjgtT5a0kuL4XMmON7XBzKfVDHHO1so9ltxlvwWrDRFzrAu/TzRI5d/QpB7Gja
gsJBozJPqhYGFZrpWFAxvwpvWrnpPjAljrl0ZLh+WUOEQZenoaeMfRldxtiJ0BY5GBtU5QfZHkUu
HjZ8D/z5J1GBiAq+T3A28DNU9ocKERB+/wCyxY3G1zvwe5l++0ea1Ht4FfPnzHQK49ZKAKEE4Wgn
aRviywWmr5mb/oKxv1HtfSA4E0ENm0yve8/cobsDIy1KU9Ymb/C/oU8sioI4vLu6tZF5xet78rJo
kbtITmmqoM7IsdSAJz2PTAU/1u2MNo7YbqcXf2Z00KALHIwZwLgDyJexGfBIQBND/TnljTcGODQ4
xLL3AX6fO6JMmrEAhAH2gRtF7AXK1zYiWAxVHCaCbkPL+yUo5WxJv1C+IZk4uKvyjFdl62QMR1VL
1KcL0wXtc/eJRfh172nV1bN6l0BA3RxH2NV06iega0TbzGrnyYEdd90VT/1gX8mT0d9uAi8G3As5
MqLWASGGh3or12K77ipfEnwLw4SyEfRWK+pi+SwfIxqIwi9Xg0wr6UkkiGL1F92Aw+NXhgnfWdMI
nqijxB4d7bn8TyhibvNYkYsdUgV6Uk43/YvAS0Qcopncmo1bY775MCVIUErVnyXVND8MwH7F7bT7
NEWQWDHPodb3OZ1cVZbtwybY/gw+EroAoatkLF0evtCfccidAJ5a3zMKzGvE/SUwis/B2HgtCYrB
uHH8fhhcHMYLCeKc2N0YIq5fu3pmcNpFLRWNCAd4e87byEK3puNfh9vGf9FlVho2ZlSrIh9iA1L2
tmDv6lxCpvSTaiIUxTfpxWfdoV6MMpJWMIfdnHqtlrZ5yGlSbLsPF6DHGp8QylRJvS10Ji2r+eRk
QHUmZ424vAqjqBlTtwG1VE0XyGy4PdPFKak/2SDe5sl4KpZCVSFdr+5FpETgmuRRSj+WmjPEgzFx
O5HlPRfRjlrqLmN6F7ujztsydDbv9Oe93g0BmUZfGp7ecZ39/P8Gd92MboIGasIKxv5YMv+YVuhz
hQswsPiEnfATNSRbi/eFhHScS1nwtDrIr6Arouawl0+jbx69DKmgDS2GELW7UKHb4IL3sCF1b5eD
t8RNne78XPSLPwtXalvq08I7q7fy5tIvAK/fAVlAtv3hca78KtHptAnmlTSm1OtG2/1ggF2shyim
OGSGppVc1+SON5L2v4cXTBGO4AQcjbPfXcwdGoBYqnyRJRYgFvz+p+OpGIinRsNuhuJmRcDQ0Mwz
sr2WRZm03IkQawdAjBS0qiA2YT9U0KujGtb9tyUT2zLHbdOvClovOnlYEQU8q7yOxO+ocDPG8tSY
STbCrh7EjTa19qEzP/eVCfZzKtplSFLXNdH2y5B0VsJE1QvyAxaeY3ij8cQNGVnEIF/vq26//UBR
3/xY+6gMqCW4aPOGqm5QKj05iyUlnyf6SeeawijULdVzRVDqRC+mE6obNlGmopcdTj3hhitmtjbW
SV/wHGM27FgOhhgCdTy/OCih8kNqGqbUQyBjTklH9eT2FMHHKFm2HYIPWoqKD9gnwihuBz+YLl2q
KkHCSD9HhRiv2812k+yniJfku7gs8bRjNsEVeZtTZyWBJZRKisj2HHYLuckWylHvy7yGNSxr4lqx
tJaipCn+1/fH+KeH042jfycVgNxqycnL2quVtDPquKhZ6ZD/lyNw3nmVGQiJdC5lfmkNA2ifVddM
xDZ4jTIMGUla8XQL+csyIM8Vv1g31AW3P66iPrgPrKrxU0Nt8BJHs1KExzEjURYL0RDavGX+xhlc
EPH7TsQBCS0FniT8MXA8PeGJoKIHiKQtn3XIWA5NQpjqJJyllC0oRHM5wLAYPweR0ehfOMGQIVfu
OcCigNVk5ukL0vsPmlPJM27Y+LGy0daq7NiRcCAvL1HBE6bvlxWz4OThRBBI52Ch/Du5bgovq81W
ip9QGALgV+nZQ4LzvKs8gI8y0GI2qKZz1GW7jl0KgRn3kBaOoHsog4kykQugmLw6aHbwR7VGJ4Vp
TJoe2nGr1UHm6/uA2U4dHguA7M5IJ3nT8w9O1xpr5HcPR7FD11KTU8488n9Uskf3W6A7LMPyMOhu
hBTC5CAZGaNXVrDUOxu80vLnVci4qOZTmIkgHLVu4JpkEiyurSSXXwnqBsqKCnCiGJP0NHabYzEX
3CrYKLYmcaJIbhqgpjqaacJkScqWUzzD3Xfqni23dHhlozIxYIBa3t7i+TJGYvq7U8X4/tpILAFP
5bfbjoicI2wLH4Ku2pBsH1ogm1YJaUsTbTsZ01+u+FJdCLdJ+pWcw291xV74qtp4GLnfVDedLvwL
p6qA44CbYBNV33dwCk7l2Z5T7MIb39qYwo3WzraGgBRdUWX7I6JxNa8tB69LVe7LvhSwmAA87jWJ
WhUG28j4fz3/TjfeZJYcTBhPogbJqt69A7WdHuPP3hNkSN4hytDFuveG0yhi5HebYCDKTHdoZ7XG
Vb5kLZWXOP0HUA7ckfikOiX7ft3BRvfVEBucCl3S6qqATiZTJqeOMjK4AJjtrITSNI3Y0O2MAGyN
PLYpA1Gr3f+QnoYqkeVIiF3ncLZrepty/fPjKCC2cHczHLMYszkw1rkAEBl0Vn8Rmv2Bl8uzSVzC
AI4iLFDFYKNgv69rLk/6rS4WYRweomcY5Batv7Ie2YjsVxbF0O41MKGRkV73UdFeV9SVMwLFNSti
j+f2Cm6qjz8ULwakN0vZDQnWOXnt1Tt5Mdoh4OP8p5CXaBK5H/wLEGVoxq+4FpFb9AaupcxDT6Zo
3ZYqAo1svTrWHYSYK8lPaqipaADklUKjzx+tNqMXaIOHVVtadV6KMrnCailSWUoR92wiDErSmqhb
LZUrs9HZ9VD/n5UohNEksrJUtPrqSiq4n5HhDZXF8lCKMhizujC3iFnGDAGzFz2qpCejLLgiY7oo
XB4RmTTLOgGQQ2xveYpd/+Iy143TT3gluYXrCKh5lax74smrH+4W06yUf5Y/7uds1cFIGRW9FMzv
tTgTkTN3FUfI0nJk9v5TpYc8GO6O1t9DmvT4/4USYEKYYmppMGzG6a+toq3RV6qkIvMDTwYex34E
c91GmRQkAuEHao9ByL6E3r4czbt9HdWa5CR3cmoBCDOFjKCB+QMX7NiQHKw4X4SQQdJkN/R9tDml
FBlSux6Zug0QYtmgyWE0pqB1OnuUTYVuG7JV+AXBBCcPzOD/g8l6mxt+Ub2Uy3chhA784rNbTM/l
Zqw/g2uZ+JVCesrOK5sbk8p6lR6vJ7HrlABUE4CVFqKQbfOolI1ogVyCLOKWeMjxHTepvb4tWym+
qcJBquu63j5cM0YuFCXQCKq/Xyxj0NT+a1mnUOsnBp3GEUBXwOlSUKV4sOtFeQK/fPatOO2tLNUz
U10FjhRRkBZzdiJ0eV3Zx15xHyz1AwTO2l6fynaVy/XXlxTtnwcTIWf47MVDZkaFOI+oVAnPeJ4r
ADr4jsBIBTPZKdkLqto+QVTLO8DnlUxL5sTZgWgzVZ2sgspGl3PYUhOHmS90TVt5cCsqK4gzXqbw
NCN4IRg9xnvZuS0xAg2fO0SkNZvHr04Oix6kgLdCBTgO9KmAjDGACkeo5A2LqkkvDRFpfE/ejKBE
F2qrpGHskuP/0UsM24rsTbAwYMeHE3iKWnsMwZgZ7pw0jlEoTVGvqWQFdRM9GRGQspLv+VmKi6Gc
RFDj8G6IkMrBBQSMWoe3pjZBgXpyxpJ562tAAktFeqyl6awUGrXQPdxShHaXrFTN1WtFhZE45L0W
OsrSQqsIdxQyzV2O9g6j3iKD/ITI9oAOvEpMcbi1r3dUgazrWWgFc/IhfVa/u7KGkhQAt46XneG8
en/g5cqYs3VgGj2AACzyWlWpoUCMO7X/90VkK5OaAzPi/Fw7xIJ60A+1UXmSd/A3l9J6gzkb5/h2
3C565XY36sq9d+7N4lMTsoM0YDNFsSqypPJh36hFzDHdOgjS+UknshAOHyyL2iE7MYa+1z+HkLvg
K275NSGpqMGiOv51yGBqsSWA65cnt+5k58CM5mVDwIZceysWE4zqaRlkiqKz5HPvC3X6MJPaXiZo
eSKMxDNvATzFxWqCAKbaICwkZYlDm/Qww3zrZXdzj4roRGh1ulSiaoIcVcuOhXbw3/f6JicvcDpm
u66GbLC7YgqO0X31Yp6deFz+LvQYY6IiAzkbsQGZvQjNQlTQFz40WnH9hmJZle3Mn/nqm90IYnKx
zOXdgZ0aavzihrj8qPGfh2/870WlJEZaOMWBPJHuokaZD2VOC9S2It6qRMCGL4AKSr7PjmZnQaVn
X84To617BVhXzjhacDcGX9Y2o/peppsnmWxLIFK04q+pZU+KbvEZeyBOXLE3ys93Cca38BpLFqW5
dSX15v310IUfAG/MyyapYZ5McdMJfp8eLI1VnzePDt1DKR4Tc6VmXHSacqUlFf9uwiFz+SCGOt6Q
YjbPqHjnTQLmqnorBPB1cFIzGCekN6TN9jBQ7J0SfrPnv4nt0KW1/tHR3nq6IihlJKdyvqvGwZEK
VCuZiPMEEw8DvWOUA7m1+6SfOGgRFp82uu56+9OhN1P+KP6YJu5BUxYyMd7PtAALJfjIQAbNkJoT
VJmNiVypgXl9iVCx0ausesgqOMlAxdatWFuZS7vzZ/pdfuJpvc5gXvgocw2fs42qk7Y/4JHJSeBm
wL8OdmGrbUHiloevjRsAnRaW4AONAyFHLRjbbXKv0UJz7uFXu+dWEJG/VqKi8ObvjaqeC5jskKBw
yr5ZfxfXWDYYv7HXqgYcbUI1juBtWVKjsA5tjQP7gRUH1CQEBOpHVhD52dRovnlqPAuacjMqAkNv
jhlEN9hAfnUHH9FcXEZaFwhYlr0h1dYncNBN/+q5O+k63I/2EbelRtuk0xt70+osOx/m47MOt6nr
su1b1oC8hPRgSX05LUFqVsfrhfsHiKFz2fAt4Xjt0bue+o5v4VP0ZCIsNbWgq9VTt5prFrR5Sxyj
JagpfORZMzKnMfquoRb98s9GlDORvdFVr6etrnfN+uCJMzxdGBB/hePli3g7EUJmxxQqee1t+HTO
dJZOdNpgDM65mdow17Ok+Hb4XdKx9mGbh/ZKwbFsjL2Hv6h4YCn9BFJhE7cClHtgCjq1eNY3vUoI
8L4WfHUoKVqxQ3eDKiKZ7nAin6qTE5qi/WV8zvqybAfZCnQlnGl5+D+SQNblSsQ3XjtNEZHxtoFL
z2GFKfMel9sF5FTR8gNI95yeY/wi8B/7FRdNfnpTi+Llmwc1mL++YFntXXykKm3ZxI5DSf/5AdnD
VYTzSORPlnj4uU4nhd5hcDOVPe4VoYrf6skGgDQAC2we+dkWR2iyi9GE2eAZERjDFDuI2we9OpLC
Kv2eRkZTShSEkycvVIlJsHcFya/6hP5kbphRRrE+ZKGN+qUGPoZQ40nEoUghlNQpCtzmJMgG2NqN
JXRWfh5BviPDxk2awYQsBgJOWrAHgKEQ0ON6ZRbpwTUgSPQV3xN2aXXoijnO4KOI5JBqhlGmxAnq
fnmmvqo/ZLUfF4WHklzOwBj9EtU7T/DIni0CyBgdQ9PwTBU1jF9QlZJJV+CCEqYYS67Xwf7ldKgi
Aw82UhtSjwmlh2skXTTGpEpY7bcY4hexa/0JeBoKpX7PZHwi+sDE2/aM5wRSIspgivaASxHU0x+4
XzwxkT5RW0eCQTZKM91NBrl65+v6U71BuQeeYj/Ti7ZlHvB0TvMZO0c0DJHBm9GVF3eyV/7RRkl/
grjkU4k8J0OTMU3GAAbRcgQ8CZ/YxMmyLQ2TJQnhrX+g3AZzi3prNP4m21U6gvWyopk6/2GdUOM3
uhmo4aLBNBOddSzFAeUA7T8dcfMOwlc0uzDGUdveOE1ZRa6iy8Vqm/IlVQRlMSrHj6NL6uhsDmcB
JBZoQVGqZPPHjjzSklDIy+VXpr0KyaGDfBpHhX0sPls5mRiM3bSZ4TGuOK1ClUyZicp8HwqGgxL6
+nF2fQcYnrgm6bU6ZVd2M8HF7CkgKwFNlBk1L/DMQxY3dj2us55FN3ZTgIhEom4mLU0Q7mZBCppb
57n8YHtRCcLRw6EKujrTzG8pt603u4+HJbNV80Lm+Uec7My40OeiyIIJqbVMhnozMD7XMVxesEWZ
zlWOTYbsTRxFZt+6drLOi8j0d+unkM232rqiyLiOa1qdaNlzGNGc12Lk4AcAI43U+BPQCbCrozNt
Lq3N7luFVv0UojS4CbET3AI3c2G2bVoCezMalsWxko77aWjoCoVFUuv22YFf+brH9YBUkLbjvhYY
Wuv7aLWnCUvSdWGotn9NHG1KZ6uEncf6s3UE/It+9Cgy+ZMQsUa9jd8QmocvnvdYhGMF/2glocsO
U9WPFC8RT+OhRiyKtlPIOhrpTqMM9iDrzqTQNxb2tB6EwO92SFflRy8Wq+1Ibp/Seuw8NfoVM6iC
SpRxLiKVHtqlmD+GtFt44epAnYLPSZACOIV2Am5T8s/yopwj6qCN50H/3EtXuSZnepdp0EIueKRl
sC33eD6nYx9+1L11o4+KYJ2Y2oRXeFQ6SwOiyB/uyfU1v5VHoaBBnQeTmiX4OfjunIUdqiKDJcO+
6pMCOUdWX/Nv/0YSLEiFG5vk/BKoYXJ+YU9ybfIJWMGlZIXBkBa+xDnlRjR7a8QlBB4abKyJY1a8
UinSMtsr/RQhuFrhZV/nbC6rfdXsJQC6Ak0lfUx+0ZIvRwwRCX+dIQO4KcXgqBbnB2QlfstEtxyA
0n+fzNsUK8VAVZaENGViA8igMiJtk2jdWikYbBvI6qPS34hZNYozSFKF7I0pf91v/JGI7jIgsqaN
ifxAZUGxh7AU3uIo7bWf/jY+YVFvMx91qxYGjQN4XLk16r51V1z/WAfFN51oTaqTUbAxDd0pFLrN
uJgKvluZiS4Hyfghis0ImTjipZ1cz+3YdPWhLvx854alBl5Sa8+FofqdgdBGe8AEC979yE0vdu13
hUDVqDCxmAt32+apPEwS/QQ/zQXJbVfyR3qJACiLhR8fkwfLnuk28HrcKJezp7AprTRvGnyYRO8B
TK9ogwaGN7iYTSbF8R4paYlak0xJ6XCUT74DfTGwE2w8MAeoflYTu2M1saHQ89011DwsUfeFefcP
F+OBNnsCQbH3T9iP1sSFrPVIfA7wRY6lkdfvG0aY4KQefUXbvxhh7Cy2J88SDtDnlE3qOihBPaon
2heuQAiANQPdZ9IR1resNi5hylzv4aJSkVjzmGRoGAk8IUWl4Zr40Zeyu4gFYJpBQVwv3j3j14wD
eH3BgULvpl5/Y1vkd/sfDBrkRNBhDpA8MIabVQz4qmPlCrg53vU+Z4L8lumB9YtXyeJejqZmyeNx
SoG4DQlq+Z5QgtPiBgxAheiLVtB/E0YlOzbaAIPGfpXMrtdWPepD8blS7z8808pGc0n5MaGzokXj
Zb36YXjU0XIHZOwx2MajmrRNpjspQ8dBVvUnlqWwBmYFS50KA3vIlDJEHjZnXN/v7txtWK85zwcZ
SHNbTFzpG6E+b2CvhpH6Pee6V3lR37XqwcwsOE5wrHnfxhn+NFnAFFczTUECubd0SOocJX2JEpne
5domGfwwJefqxHb6r7C1OyZEOHU0f7HeRMgL9eoq78NSMvnWPCq6au1bJe3afoTyS962/JMu97Lh
RQbCSKHM6Fdk7M3nC2bxXuLol/ciTLViwDvjVkGpzzhUKrfG7xu1bRqhumYPYDCm65nzX13cNOZG
gsmNBhYNErnwYCdbxRGyh79sXU2GOp0bUFTqUKXnfUFWt5RpskEEsfUC58pb7fdLgbnFa8kk3CtZ
mCoqM/6yQL/iRd+gIp1SPDB9iQrP1qP4JCpIs4BvB/jYtAuC67UvrIjUiWQpFHNVNJxjNzQtDWV1
W6r6frCsBHH81LqM7wcscSEIjxYW7HfDYXA6q4BtpnNl0bMNRU/LZfCOrv477A1FQgm+KikOTwIa
Bd/H+sN6S5jfAmkFsj6uSnMCVvUo9PnMo5kNX1A1GvXnJBZ3TK+T+uF+ZNItGvx4pq00+gor96lx
slYuD4JccRfcuvf9EpXdZHyU7HWAnCUDeTJtZegTf4cY2jwIPL05yuBPLhH/UiCYy95TVrxdZ6GN
2ZBlQDuSKJ5nLLGfaMXU3kOp0lGEjWpJB2qWL/VDeH9Azj06HuliV3yd14g+j7as3QiklKPmTvzm
N7uZvOK0nxIXbAiGfdk9+u0eiJa24unl4FlhCgxH2baaa3cr+U/Ay2QS+E1fOYjAtUyaahDkhNbC
9oYkaG/c7wYvh6zWcUrHmO7TA/RDdd5/P9rbe8DH9RxZkKD6eTYCCxKFTQWTlNjQ12ljYnyU5lBa
GnM317acucQA+YRUA4m6CQcWXErTw4Js9XeB1WGOlE3TtO7okGQ8LTKBFl/UJI5rHGOG2+0yrw8n
BSq2xHOlcGP1ryz+6JIxjt41tcSH9KChkjkKYOT7AVhgtna2WYVnlaOvM85xt38Dx+ftGAc/T9Ps
GgDLBbQNTb1Dx5xB22Sw9A+C4B4V5jDJI25tLiH4Hufk0TRnylY6Eo2DLh/CZRQZ7ZVunxmTHr5E
P3PdQzIFMCsfmAhZuHMVTZ3YH8quYZsQkvQT1lIm2IFh7fJEC+vfH4Ou9Ai6cvVXe/U7itIJ6a9z
GnxA59kwJEkK3OAqzKHK7nlmqhrcRtSlvt4H641QwBWSo8VhnNoEMy/L/p6A43fBFYHC9zj9sUMD
O4BPgIV01ikNuzL6EFSdfQBJpWfZfVx/TmNCRD4FedZdcN9RgmIFOn8txljRX7QHo+R4EYaYFXyG
ADUZCjyrmR+htIEG2KbEzVm9jYS0rE8JGm/E/6xzave1VyHxY0vwTov2fXCy+w00XWMJdTe4hyB4
r27Dggwa9+aWclGy2jNwRsqxVkgYb20ai18NzI3WVrvmEP+JqgGQL00w/qGVjAUvtCWhgsxIqhV2
YVblT0qTp0s+iacA+nGxCe2qdjWRsXFXYA6oJJOgxfVYBZbCYc5iFkObWtZN+i7GDbjzuUxT1z/r
0yy10Ng4Owl1cVP/xef6KG/JCdrj8vjigtv/yirTHwGpM/ZtmsHfNMEG3v2n6mAom8J32GFDLWYy
RQ4UhSAVUL1emvezNEwiLZKxqTg4zOGWwPpZQ/J5v0Uk6vC8GhrHE3gLjZBq1BPeOmhSSgZC42fc
75CYpbQX8DRPrTPLv4EhRlH6zMbEdjfKwHCphncSxcjAInGd1mqwSQ8b6MuAFWR28lrtyw9Yxvtq
TMV8ERa3hL5wT++zEh8k+JtxCJSWIWwjzg2zE3/A/+ay069BVQrnGWQi1JHXZRSGOMN7YAA72kSX
SPvB1LYwJenXL5vKpnBTtpQeLnwPhcsqvzMAPMqgFwJEQOQ2o6J8BXGDUeYOnwcWp406mWu9XaBW
C80kc7IccL8at2XBsv28zCXMBsNJjNznfI87RBrs/OJLpWJ7xdnIl+o9/RZrDISBcVU4H3LICf7g
5Wkjm2kkPkRQrMhCgTQt8wpK50M+gVOJ060C82BN3YlQRRkXWkIhe+/c/9fwGy+AIyrbG1FzCJVd
E69HPaoN6QAqzR9+/MplOETbIBE4m0Nrcub33RLVtOtI4elBX+jSUoP+myf57b1I62QD5zr59ZbD
J4MX4PiIn9AnB4KziUIzZPSEBt59CJYEEUBZHsOLzJVhdilB6EjQRL2An01pgjivW7RjZwmSEzyt
o2NgHfEW0jtmsaPBWK73mO5r7S9P8Q9t+EwElaczPpPqqeXevjwRnzo/aMrvAAfEQnS8HOsavQkx
iw2fY25nBMrMQAmhA7hiUjbWyLhaksdp7zn3f2VDTfnGd9nmL9FFcjQU51kjL1Bcz8/KWbHAENJc
FDOQW3bDT9/g1UdTY+SciFAipl3xJOlWvMExyCT6TAU+S0PpmAaZunLMkPXfrHH+OPF0lKcIZEh5
OWGqfTTG1teXSXfSO9abWKOAETt0rhKFxqPUK+DDDuZmpHqRzzLrs39FVWHzSquydHeCUVEHu12n
kxSq3n8C2mS27n4mjVGgqJ1Qi2FehJ+CU5q8cKAoXEYO/hu5Y9o2xJjqbpOa1CXXNMEpEpEfdDHD
j3cJ+mt1g+AD8kf1YJVvMhDtWgLt0crQWAWif0iAkcoWW3bCzp1NgVXL8yKFpxSsId/VhBhpz6DF
3EaFt2RQlS57hlwZSpB2EFBKrOPO7lBR1EMrUOi0vJbXzqRz0xGeLGOti8/Ky0lPExDtNwJ7aOoe
2nke/4PkPtDaYJ0dfHUpwP0HE4/OuViWpE87Lh8sN4SS1wjN7T/80xJSygLpjq1RlWuNjVwwOLpR
6whTkUd2Y/eLGiDumpq7xKfp5ZeloHjX4FLH0T/SSQiS515AhYCWRXv/ZRJ35HyLpgqPQxILjgRq
3hTfsDmn0d7RrUMS+eUYDUzxMUzKodJdvaN1UNC5rOPulQ1Xv7iEq0WdJ2aTJjJ2rMywQxNzSN5z
N2Htj24WPmzNjUVb8HZJ6K38fjg5u0TqCmjhCuGuhWoyrRDfbvwiyoeKRtFS3eqimy3pudaKosPq
1CelMid9x4uq0wQHjP93fNeOPY1aWCtLEQvF5p9p7nrKigS9yghf2ArgaJBOwSDK+6SYOORpLz3k
KvsV5FgtHzeMXq2T4IMDqWs7FrABOWtUvtUiajSJoCFkfHC78XvkL63xFCO71YUfKH69y9/Y7nYa
ifJyEJNakkv66QAXbaVEqZZa7M88jVd6ACAzQkxKbx3zpYvJ6cFXhdelwkVT8OvMZN1bpxdAw/kQ
NfetK34gnlz4RgUxOKDL0OLdyTB0vNC+cz91XyxaCTkjOyMCLBl/pQxtSPrj+i9fP01WoFOZmO7n
pemwuSWeQa4onXOmeIc9JAksBOQMCW7qU3yJ8GGWPEPIO0y5ePmCn0i1d0tQCtpR24LKmtJnh6sG
IBUvR/qb+hVE77jappcditGjuLLQ+hIdAp+zEie2S2K6NVeeh/SEShSXWYKNFesd4X36l6owlkmc
EDEXWFTo1kbEY++HMwVQ77F0qmTUB9UsEXCqg+Xb8/z+o0Ne49xZQbkBYK0xRbw2/bdpSq08lVmo
QA/YUQppx5KzWXvBnAF/9CFkXS655VQIrPAWxccg2Wy8D8nEs364Jbz12T7419fgafuVKiYOChsg
pfsSloClqEaKIXKwpTdM7et0U7Tmk3bE/trtVp8y1+U5akJlLCuzeWDhDWDVWe4b99SwDdrQZcIG
p4MdvVrVjeYSnxwbHODZPk+bLqj2aytKRcbDHI2CbdWjTEZAVG+7BKtoQy7Gl1g5Z7VudZC6+n9C
YySu5uR22xk4hD6yZKJeTfRCrrE+bfKVaj5X2UFhFCRZ+/DDrM27axcEj+OELR8E+ZJ0wRDXiqNO
Gkg5gZLlu42Oi9KN8uy5zKd+PXgxqKH2Z5XWU5yEOeNM9o18MRWwKkZ42JMbpoMMtUxT9UPLbNUm
LIeYCdjLUpT6SZZjeo2AHdt8BxuprEGdW+5qVMM1+FuIJZj2+m+9s2aeALfdTNvQsGeuIXjWZDu0
rp1WqJYb+glEgqO5hFJxatQEFCgo7lI7pxB1ZOyb4pBXSKlRzgAmGLBc/ZTDB4t2hYfkOtLzDfGj
z3gfXtBvQKLdXHUtzV+mc8oSThG+dMVYFeSJc3gVB83mc1mPces69tgv5j6JBLDBISX+lqLthV8r
jHkJ3gRHZLBCprN3mU5XmHGjpWaxMO3rveUw6lAt+utWv22PDAb8HntqFBBrW7SpOKAXgrbSnw7L
SsAF3GgrLOUdyCO0fNMp1VEndPFGyPUcRMjcGy1OAsoG2RhGR1S55DjklnNa+MDpx5Wwaz4LADMY
IMYA6WAjDkYBfttxLEWco7CeDefYzjmING8N1LugHsO9ZG9YpMsivA/f76eyvoGTCgYG1lwq7Y/J
QENMP+sV+AJOklZTDpM6yUugpTgiSXDSMTtST8pJHfEimsJBeRVNaTj6R/EtXiGlPH9M7QrKJW1k
lYtd9tRzU2yuO0jkCGf512D3vMVwDwnoP84yaMfOixCN5EkP8yCNtfAhuueU/a8JNlz0DuHZ78fB
bmCKXzb8INOWkDZ+JDS7kovdz/CgAEIQo+skrWRG81bJwDLF+MJ1fjLi8ic8sEjd/+nJq+lcnDgG
O/OtbHK+rIkX1ShIkfXQ9B7xricR2KbZRPcqXdjntj0+QidHJnKOAn+zF8s/T+wPn4U56qbxV86a
Ht6cRGItlIvxgTJyTET5yBzBPmZy8kjp6LuUX5UKoqx+YYrkmFSVM6+5qe1QoIrOIUbC/vPPjW+M
D1V44QF/KxSyGQRbv5FKsfhaGPDbYnKzTDVnSujJ7HT42bo6TSjdBn/VNzNQlUoVzaPhqXwNpSgJ
3DLRcu4MWDK9QHgBQSYgqcJWQNDHMVFKpH6I3RFIDXt0DBc5dMNUI84PCDxRF2Bl+HBC3Rlk3LPP
7VHIw1z3CZJEoMrmAtdqpMAlNGOLYFMfRkpcOlUfAbrC8BDRWfVe4Bjy0jYo1gHNhiON8Eq0ZV1a
U+zn9SpUE9lKjuKrYaC7i8EjIwCL5SZl00TM3FLE7HFBEZP9Q2ITqU3/+1q7KFpeDPm9YYFKHmMa
FqB0l84CBWq0nsfabbIfiNldpIvYYnr94nmKyxKVCYavbioYQX4JUWdRKMVyOIaMOyqXTo/lxB0W
YvC5xXM/E2ZuOVP6W/JKibwfegzooq0oVlzoYzmsq2K5unts3t++GSublqJFM4ZNbWxechBHnRwy
tqR/4Xfq6CqWVpTcrfQbMb1xMyzLV9RRtoblPQsl03DeYgwy4XPkfWCFjDyD5AhlAQfTzwp/rqae
R6Hl+zNipX82/TRb63OuK7riEQLaIBrJXCtxScnZqUDS2vtXEWIKWdCJ+Xhuw9j5IOz7Wx7Bzd91
65AUqLEX6ejZLxKa70ip8XC97FvDMFL7ba9aDnFpseAI+iiw9s7Do/iPjxLQjyOlAO8/wWg1pOSt
7hPZxBwrFbFJWPHGtOaIxZHXxBPvj4k8BMCVSyv6yLRwZHH9iMr46LX0EvqAVpnjJDsYM01vLcQl
w650QStrz9ZPbV0xjkE4HWse8d19hGlXXgHwhNzj0K/pznJYmV5v/Gcm0AQtfgMw9B5tKL5DVvkr
1UIv2325kdhjlIXi6xx9Z/twi4SmKjVLMx8rtQRIML73qzzJA+WcH45fIQiuYc7TR1TiqNkNeCZO
/UWB/SjXHIxlaKzuYndi4GeJBUfU6JLQqXLG5TeVCfEVi6uRXf7Qe5NLNZtTea79aua8Jwb/oSv1
/vsUEJevFsfr5esjDTs+4axlgKcQr/dR2v31eTI1p6nhrlvOitNXMmGOZnrjPiduPZxShVTQT07L
WWem0NmHBTtm5YhNZ6GtCg8EIckkQo+qIbNfL3caqiBaTMsUFM2jMKmVXp2HECXTqsZELpcUJ5V5
ikmEysVYalZPQMUBfUTTyW23Jh9AUpQ74n4DT5Iin1n1b9sJqx7/SQ38H5VFVe9O77biD8Ip/jN1
Ld63EmxLMu4jFTEtP5g5qY+uQ/8sxGm+ki3Td1p7gxHZBh/veM+FuSV3J2q93zsBJb5h3fssjRUJ
GvhKfbfes4gazzE/B2Arpsavd/5RAapwRPCIFRQSkgRBxtUbanCdNuGQid9kUhPcXWJaYQ+bfcjj
qepEvQqWQJ3H0s7AmWX2AQDCDCFfmYqm3lovPBlfGqhcCiwdbUCJb3fIEVEeMdfM5mELcP2Pao5F
q9ZGB8jacZuDzeHEYw+Miwm++7OejlhkZMVM0zUbSP/OwBbXQXiQvLzmfPmujSf/zXRYPtioI5mL
bV8lJ71Dtw1CPj/Bi3XridwfFIIfXX4Pcw1r7un1VQdq1v7U0sJ/Rx8qP8AVTkjsIoPciHc+d7e5
OEEsY0IRgVSqyZJpKSeCR84XKjfyqm/IUAiT+KnOMGA4+QTMlcaELGMpe696B7J6N5aDd0TkcdB6
aQ6zCreWhAgxa3IWMUK3FHcyWHp2Yi5VlZlaee/kGsd3rFS7v+s9+2xeCers38wP5saYovQPAf3l
HD4s8Z9RIgIuyadIFRTTdoIVhB6NjTQcznFIcemIQPp7Qn+6X3blnyXfNAcmPiP4pD/K7bRl7Et/
Zf1kPuXpZcsbo539uiLmap7D68yQGctDiIGhMl52278c02vcc+xNXl9KEbVuK8ZbukXfzxzLmdns
3su1NjbUyHtrrEPqjg/gbqnNMo8RnGFr1SNkR4AlJ+Vx+xPYmM8kIHvpo3TT0CUHNW0se2D9QTQq
kdEaMm7h53KUtNr2EtK6WhpoZmjObkJvEvbnoH9sNV4xs6LlJG8yqKlNfYJ4x+a7O4e6A4qXGgH8
6HI7TfWD/XXe/qP+PVUyS6nm+WSpspZidky7zky15FPnNP+1pwTjdmvOHngqh9dzbO0AJ94P3mPx
r0+FpAnoGbOnrsJR2PKyixBvSqf7hBg86rJWIbDjyA63MZh3Xp1rwE1mzeC/QkibY0YMYgyYmgzA
CuFE+M6A2qVofF+jXPcmOoS+7QJas15Hj8lp7H5mpVv4JlvgqJgZURzEkUNH+7B/V4bvfqeAN7QF
U0l7me0XZorboLZ6NPIDRiqKXmtDAc8H+meeiYZ9ktjZLsvGbye/JzBnWTsgFkIttdQLvpDeyn5Y
ZgGUclGejrqcmWx+ILG4NqVv4a4OFjAb50JFS/ZlTbkaUFQzTcn/qYjpLc05p0sdcZm3RUj5BNRa
UZ2mD80sJxv4nGDz4UCNY2hMW4q7YNetUZr48JNdMSk5ng3E+CEjtmDAQ60VX/ZPQszJ8ASdZh4O
Kmnmx+uyXGi+5kyVA4Nbf9xMSzwqJwvIr4M3vym9MVgqyqYL+Q7mi7Rs7fSSoK16M6GdTWk06YZW
+1nN2nohTbnt9dS+hk0C14SaDa0Ue+fzHQDkx3ST0Hzzqg4uy2iB6FsFhZKROXXgdTZB+JlXzWdU
Ov6dQUYEvc1MuDuL2Cum5EwfywONB02tfnaUMc2H1qInDUq9DKl3VOsTqp+9QdyIBGZ1vuEiR/2E
EfB5rw5YWHBHnO0x+3KKx/aAwmuBzYtqW7R1NrkO4rzqnodeYBYecSx96gBGne0ZwZVkC2R0UhDG
pMVnKz2Eu81Ht7z36z5BfrOBeKX2z50GWviF39huvmkmI9Fb5Kewu4V0bIfbyap0SAm26nklDRoI
+x6Cxs2UNbz+1gDRcoDdp3VEdHsXJctzyM19F2NSJ7hOyM5I35eRQsca/YjdF2LvmZ+GKIgvC+4t
pAfGdpApX8h1S9jbXfgWklEAonkgAd7NP9FpnGZDUeKRwBcQh8bzodlVp3QoeGsQ4+5w/Ood3tRu
wTZjcDSxOxnoXSi0H20z6+VwbvyLDGV02m/K0W/p1y8nwqecUKHIws8jgr9q2iP3RMKlMMOh7KwJ
pf2appw5se+O4NlYOD/RJBcwrkxV8bia7ZzNXKUA4gpCSCCC7JXdrKRFJOPelIA4vhltul3EIyef
7ROOvsrJA9p4gObT6IKY+6Gl+GNlhU900H1qTmyYES8oEEs8wlgidzxNBq/3fDV9sx/w1M9RwOhv
zsUiDdiUrphfT8YHOSHd7ZkwYBBclQCLm1tHZoM2QrM57L71P76fthRzFHEOM3Sx10n9MDUmotLV
Xf7iYEV/jKwRQANmrUmnaQi2iIwoXtBoR84hpIYylU7J2WmYmvf95lNLggBZNK5z2xp3CuzDCaFB
IXF7CJx7LvYZXeXk4bHXymY8RFpDyi3D4HRSlJfEhbtjzcxGcrU0fxFzfervOoWJSdyiBWQ1HNvL
eHTeKLmdSQMPiqqalqSsKR4VPxIyd4JMoyotFFvFIk5gzGd+qdepiANfagoFa8g/C0vXFksVmyO8
qlxnFruAHy8dzrkn/ZmXy77wk7vS1QSOIZtFb9pO9vcP42ywKWpWK0/thLTS3SXvuK/bZJIZaZ+2
VFexEs61mJUTy627ootoQEKDF+h5w71MMSax53jsbrRDChRuTrbpqhdjqP0fEOt/5H+KAGQVfyjG
Ul38pUF7wQWWYfPx/HQZe4Y3p54zpoQsaURRI+VHaozekb3+9XBrsyn4gBAt0Sturd5PQVPmLd34
fJLQpijLYNFklqf3/bH5ZIC1UjPBGBIg24RkhBG3QTLsj9vjTVb41FhzJvgKdl5II17O+t3h+9uW
5Q0JXCJcOV/2qbKOjFRc99vjEnX3fO8M3+LuEZbcCfc3ymKsBss6eVBbO8lBKiVpZrkJpOx8TQUr
s54bPWkyN3U8iKgbi/FGaISq/Pyma0cqJB/s+pJ1l8DQdnIxapNs59EO4jV1ANG2cIcO8ubfXgF+
LsOqTMUyB3PSbovi4Lb0YoO3bp+7XSOYzAnaXtpTNVTN294k3XmcynnyRvmMbQBUEc2jCz9g5bAZ
ripC8+JQ1NJQtHE1IUS7X8lfjBdQvaofHeEiV3fhpWIb2oKsfmpIDB/DVlUDQSulOA9/VDdZkgl5
+1GTMSIKl89EXVE3Isj5n8F8nnreHjb36N9ztGnK6tfSjFC4FvLHxjNRrqEss8EXcLo/sfdnUPOD
W6j5jWC7qQugrxtTCjNKUk+BCy2lA9tVfUOek8WLeEp51k09XqibHkeBEIFRoVirdG/MTvFeUMYv
WrehzdJAjMjHpc9dSpFgTm25pbK9NVuXETQebFaN83z5IMl8gRhgIC0LryTeSVYpvgIQWPbkL+Ek
Gxkov6wCUJTKXPTvZrBSZMA4f87ZX8rlumhklpkLds9JqbyWSWtQCSIDeQ0Ek2DKkBx0Dk3vh61R
Xg0fT+zzMRyB9TMj44MzUIURiXcQIHI/oLGLnIjqOkrk+4TJFFCtbmLL4ylWJSE9qeOWYgCleOBu
kDJISUlG8/IwFggSFFupt7pNdAUZb65Xotx5bOXZrdiHARTU5p1+rg8lEJnorn9e/mC/iZ0And0/
0EcPDLWh7B3njajWGKgpr7PrHw/r2l3QZ1vDA/SnwLoBynAKETl0k7HAZARd1+jWy641dcDjXlbF
ssoHl8RSZfB0nkdX+paZzOwxzO58nkwrUrRSI5u67E+iWB8qovt1JtDwThj/t+ZOyhmOs7h9uVaL
aFyzL6C+33mVr8II6YZ3b3lCGFRRikjQl5NBpqWrFhg++GZVpRBZej5Q+DxvA86v/47M5PTFJR4Q
0wgkFpL7PzY+xJ2Ete8Q25OYx9Etg9YcAgxt9QWkxZJ9pRNT4dsIF4hDZh8lTzs3RaBOecVGwMKx
Td2/D11cFreQeutrwpdhpuh4hD/P2hwdzcm5YnW9b2Kc3sNLr8pJ8UCriWTYlnGTDjze6Aelwd4s
6E8GAZkFLv96zUDf2gX+QZoDILBFooEXCXB6EiBr/RrgUExm41vVwsAUQlkQiGjJkDaki1KUmUfv
lfMt9wC0COGtzWa+eIQeiRpX4/QG0LBzJChwOkWwl32g7EyT478lEbbNQxtt/APVai0TRTcg4RDB
qbEVq1NTruTEbJRn1OOqhh6b7Pqgbr7PLn0F85GJSmWpbaFFe74Ozq+q5USwsYXmMpzo3kzUe3HO
Maj5K5q/ont3yORQz1yamSjC7UtitfNlvg8gZvXQUjUMvHNgKZR8DDm92rnKiY7KCIdJAbnDoiCZ
KwPK7O3otSA2COv96Lae57l5JitX8eFtp+V0EhakYCu63TRc8OD+BHvLqVboUtPWzOJ95lO+AbQ7
aT61K24bWyPer3OzYqf0wEx271CzRwWKPRiqfBnNjRemBWmg1xcf+lzY+9LYKdSm6Tjt1mXA46En
p9lqPAua/n/v9eXfEIix9rDWbsarA/gLU4UWIXddBQDMzh6/S0qY8L66eq1crZexSiG/eB4fCqig
xSCPkKug5QE1VlGU7TRvPx3Iq3Y36843qzFbvYzQ3kGdNZis14YLFvY/+8YQGI3LkrJMv3tC3Tj1
rQDHSiLwUPHe7yBNw4TDamhPN17clVLqZD9gko6a6/2VoTYP8PvcjmFJgE5N4I4fKFnMGxP26cmg
zpCLmxK++SSg86Q4Udf6sb4NUGtxBZNRHhrwEvuAuYaG/n+5H91BErSV78nwbzi1sRtpq7JsdXEr
7MExAHSomU9e66zDqKNTqlL/v5o0h6U6xdlcQQk+mAUYDp/4PqAsbA5dqaNFN/KHX+lar4gmPUJ1
jPdfIve5CS4kqT6WOfC66VVoa+Nh4UHI+dbpQS4veZBj0lBeZsByuB+k1/2MZfgWIy5INwpS69XM
Yr3NYlU/gfi3af55avmU4LY3oe9Y+G2Mz1K5f1vOb3r7UzEzZbMqz79vhIvCVOy4LxYkXMUuW9D2
o5kp+2fs0LKzSxvhQxmmy1nLLZYiKsNBOXCbR1T8B0RFKjHEHfhb5yKlieI2xvs+ZPEIpyFUdS63
SNQAkJcv43FR+ygkFAhSaEKpAfy7xu7bsUF05IpJKOCTy1FXgBoXIdo3e1O11hnh9yDpFQ0iPOCd
wa/Da+vv687aU7lfKuRYP0fy+J3lLINrRYCV8s6/KO4+iL8F7GUGLfCnXgYzMi34poGan7xOu8gZ
Gzyi5UProRjYagBEDnYSAABs9qyLMWejj/ywWIkegwhJN6K5AboiNB2l6SeXiAG1q4CFOwQvsaS0
nBuXQaT0Qds9EVRZwnpICj/+2O/ZzWMFN15BjdljReNYzYAx3aUsH0YQRY3rF3zg+0x5/arlwRQh
m/WXRSGoG8jivy94EhqXLUSi/4tyFzwbUPuVKwPfFBdVSoBY+XajOPGucPidipveUSCgTT0V7TvO
uuqoG/DlVG5QQLrX2o1vil7lUJJidZoB6z9NwxPMSSgurw3AbfMz9J9b+IdvODT2DEhZy6Srxa3c
hWWA9TQ1KAv6oXbOGYa7CcsAC8zM+0jDI0Sud3vbaZlHfuoUzRAoH+uQq0mLrdjsED+rerUe6ir0
UPj3nkCZEmYyiK8E+DFp5iWQYkunx9aK4KyhTKzeDFXWNiPkkhzoyBpYKNZQ/+A3vwzOnEBKhl3B
kohoBsT+PzUwCqjqnZwNos3hJ5QZAOXMskHJGQCJbvDwVvSzvD9QnK5Uts32jhOQSzQqDzacK/tw
GbfVr8NZ8v5tP5SXi194LUSwFh/BtxWNgxWMDPC3ekOAtdVirBfmqmh9Mo7d6De+zP3AKlBj8lsI
mRkMOfICxXqTtLL/+wNT0L/ljCvh/LiL7VvSVTBgPQgg212j8srN/VNYPfdTPEhy49jSe8Lrv2ji
itQdZSdEtooNzbDEOdo3eeaCqWmZJNN3XLSOiFt1s4ZkZzJ2rH9O93E6cdkeNesmQCU00i8lxvwE
E68kDkGfGkcc9keux6v7w970CeOWu2Uc7/7fbe+jg1dk7437/w633G0DCVfISplkVyFhEh5aJPvJ
P5N51HuJLC8i1mtcyoMfnDn7glLPmOlSVWqB6jnM3/hwfaFAZkdzxCFQIlH6FpKMkcTK0+M9893l
XWmOX/H5MEuf5w0yQN5hWew9xt1I0YulCClqB+F2MLi6X3RoSy4oTjGPYeSu5lkyp/1/XKTin+AK
XvPm1iTKPUgr1eaLHgTtieQbzCho0aZ+hO38dZzVMduJDmCMzMcoWsfSIqfnNdEvd1llocSzhkSb
3xp6z8/wu2p5lKh5i6f/b9kJlBF30CPTc+oxCC+ZbeEXdudRe49lIL9Tfjag6+PbUlLhkjrPpXnL
jouq4cL/ShXJuT7w1Bu4Zw4mqJRdJ0fU+a/WoVrg6OwxUKZz6Ur7q/k/8vFLFlOkZy+L/X6QLkul
QlZxsp3jSz9EosZxa0+TVh+hvJsU7BZSputeV5+D+XT3PDmHkwm1KR8ai08FWUNo5Xcdoqny7HFC
UPk09x/sdwrAXIdvMirhjJWJS0sda134GDY5URsOCtuGyIaWmVuKVTRInkQbToU2TuzrU+aC507I
jG74MVGogHIjndvWi8o+1666CtPZ+keUFUwagXk3vzXC+uN3vZKg4qLLW4d64Ip72p0xp49YrZb9
aVzw////SfqG5c/NjRyZJRHG0XBxgeJ8qkAcNe8MpS7r6mkTsGutR5Q6XRkQ3/4PHJBBfhphlEYj
23p2W+WWDHHUczVkA7T5j4uwqwoQU67JpvTiD2aibrQoOwzM4nDKCto5orAlf23PYP1Pq3M7Mm8t
WPN3/SlknVv0DoIVQ54GnL20DNG4Es691AZDOGm1PJBJ+l7V11lYUs4eNpklzvjhbrARkp6IKcH3
sUmqLyzmsj8B0dj4Rxgk/VTNghSUOOl2T7vISBQX5HvxKN72GqNkcBussyYF/3ha1Q4k2CA6yT5r
UPkuMVGoCa/AVnA1UAc+KtW8EtcXNeGRnnc7nOGQpt+d+CJUI9Xvzov+mwlREzFK6nLhHWzSsLEQ
UEXIRYeIdDbL2EKOjVV3HiWT+58TdGwAiHTnujKhL834V19awYgcPfbc5mqmq1q1cBXUCJ71pNMi
8jruWw4xqJAhgSZeLOdwFSNAffL0yyX0h5RUSNNoUXGJ/gYjcYfizyZ5EZnA8UCmFTz7OYQ79Qwc
MQtg3Ml3/7eVsTpaLxZook4nWpVEQkA1yPvCpW8mfOs8vA8DvIlz/ziNlyGg6mtOObzvRIxV3Mwt
YyVm6X9JRPYoPIztkT6LCq6oYP9ZZSP6MxBmoa9Q0yVMXZ9JOzfIUsT09Jzb/UsH4f8MYDzwc0wq
QSDy2RBo+ASzWdibfoLilvbASMPjXZV16wyBDSf0K6ZG939SPYHsc3ckdYib7JZrQBAa8sDr+ZZz
eLPvaPu/YpI/OkZwyDYJuzZlHxjZJD0oswCIAfwp8MloY4prrjQM96ea30ppGK7ZKAcSxEnrYSKA
1+ZhlZUrx7T5JbyGwV9+Hu1jqnrjQYaXj2hwPS7oEbeHlzx2G5IWtklSIVIbdpVN0PXM7IWXSpeq
8KxAUZdPRKZmum+IsxYVeEqg43hRa2HFYqjPObQQQQjnZKkS6dsBFW0r1W/ntCzGwNpZaePvNSq8
6h3h5sVM4tjFmolqt+4ed6VIqHRKzY9o8DQWwBaxu0alBmWz7KPhcco3xLQ7nXZCxqA4xmMndfJd
ObD/7ZcoYDz8qLfx2dyjM9FyJXhDTf6IVMnUXOYGKUIrrG/thwovQaQqkpIgC9uEb4ms028QMSha
6SP6aprJ9oJRqIYWeBXvoI9MM3mNPYHDWKmPlCP3AUZ3OYiPOIRVnwErJBCbZIRfnvV0S4dnWH58
lhDTfJOEksoipiivKy0G+aUXcJlscpJEsajDEHJl5p3pm3XsplTQTF5BUX7VeOM3gLDvmKmLoNYL
qL3PFoZhtu0QXj22V3UniWF+JOmcA+JvqK0+lAYSndXJaKKjUsixBiBBItAFQXudajumhdsWjSK+
deB4CjhRh9aMnACk8g+KLbg5KugBBJ7U74Esmh4vOYwqyf0iZ2gJqsPhqV7HiwcpuEwk2ZRcVVGe
CeemLfDMBljFh0QRPJMxiNA4nXwAifGUGfIW/6M1wdXst3XmgWM4Kpec5tTE8j3Q5m/Tjy/z3a0X
0nm1NbnX5dbzeV68AcQoHdugbZGcuocxJWVxYpUVEzQ5NLZsMx4ozmHAzLHKx0U1d7KBwz6k6yVR
WGmUKRty4HyyNn0JCNU6JByVywDfo46FTK8d4MzqryTtSOAtOAtuvnhiRSIXOZxrtZDjger+73Uu
xoDZcFHmLIYRc864uGNOkQQK1RPak3u3f6J1pR5LJQhl6MbKrkIe1lz2tvP0mXMwvrVHyr/l9NsO
Q9k1Byser/rP+hxvW4/2deKP9wGk2BvEuPFKUJ8nZdk6mKnjy7Oh7UwVEBbkACUdyiQt5kKsncIV
0D0ABUpPe7gyw4YI425ZqEPb3iJ5GY0Q8DoSKXRdTaFhaw0pDs+/yMPX/u07EZtB5TtaJlOah1Jq
gNrzBI0j+hKkj/6lbXABghjb9dfVz5RuhgQW4zYzOXoytxIBZvrf9GNTdXpY+VXTpjvyPd9bSTca
htMVQscTEnn8RPMWb9y5zptwLlCjFE5z8RwenN+ZQKzg9NyqB49NEw72QG/erp0vnv8TQLlIHJR/
bC6m4iZBeGlUmr+R2wHGUqvdEHMbqvClpwWv8edFYT+6zxkLiZ2x4am5IR8uyZ/iO4JhltZ1qQlx
dje6D9/ltTyZl8Z/8Xr1SAz42PXZDJMI0d0xviz+8GdFa43JyQe6LaYLPBVpy8Zj50SORM91vz2v
SMBI7lyc1dtbUfwhxVJZdkdwOx1U3Bqh2KBThw0xFJA//NmpuWPLZadWi66IveN/Xco256Ghcbwu
cS3j0NA8bbmVYzQTW80rL2gBJoCeiH1sMcVTf5RyRjUJtlVRbgw6ykjIbPpbKNGhDsX9Jn1A1y9p
EDKpHyj6rd90Ay0r6OUxOeu/fY/wH9jrbzoNSAr11hoRhHPOuSw1vBpAq0iocDeDoybrfKZQT0ZL
FGOHgzd3kwyjZs8HDhTWcysfZgtAaqJ4IsDLRlfoU9lQ1vlLYasDWrbKkUhtyAkREZ4OAipm4ttG
nP5sY6drMg1GIoOyR5KXVg4uQzGB42dDCxN6vZBUJYGRYn1Q83pMfpL+6nXAOWkS3a6TcOGlBRbR
LVRoCnSR9zzYR4DcbNvVbHimGEB2lQI3d5+N83oP9NHTrjBe114czI89O7orxrBLetPb967X8A3R
sytrkSHykUCBvOcb95LEWs/cjc2P4Sk6TEM2i82JP46Uj7WfcHRkgJ/Cyh9Of1dgIGbQWbhBtQsR
dwDSaDa2W9aGrsL8sz5BfXWzcnIwg885jQ7BV5GLtln7/cKCL7kpmZk/H31n3wl5rt5P3b+C3UDA
5ZFAoSvwQYshhtw5sta2jXFYkzo4UsJ+YD2bt5vYVIcbbVAw3TCRQnxFXXrVKX8h2MsYXvJj3E/I
g34EIw3tLFPxHDuGmyUn9bEGQbsoigNm9mUTadYV1auTFichfsfjoZb1Qh+uhKwDzoHWsCarjCJm
38hJ22JTsM8XhNnJuYAdPICzk34D/4NJYrDHr2R3Rsyd+JXzLMAiKo16fg9XNaURvXQB9KFq1xIk
7089dqZDd6ev4cVKCUwaMAOLLXywZTXN+8zaJZxGUCyne54maa6phsf3mg/R7U9VjkFXgLWa4IEW
G+GCT8M9e3mPQHmyWmdpvqBC7ncKU7vIt6uFbKLqwcy0qLSBRE1ulkgcyDms4ANk2s/HC4yAzkPw
9A9lqKUCyPYqcG9xK0tcyErpP1KUPk0wrQc04jdX6p1tiluulkAh5Q+ux8J3c6AeYXGEmmOc5gB6
WJrOjHJusemWXm0fE7nmctXwJZ560WFFcTywzNjT6R8hd8VdsjNSePq0D56X32f/z/rbKD7q3xsh
wkR8mbZP3/Kgwkr8Vy5eI8D9aB+e8VZ8bhYFB2ExYaMtEtGqKl7Gmxkkhi5KFJVT3aLV4sYjueYe
IFT/jzVdKEPgQljgHfcJ7lJifmyhbGFwhYdldzcVWtXBWHzfPBju+WI1Rx+pJNO8EvTTHO65UAnB
W9OdjYxlJO/QMax5jmA9LJF5yyTn56Wk1cgaebLv5I+3OTmJk2Qak/sS0oNeTwWTNIFiCZzrQpAm
1wOe3uY8MHbJV8kptwTqywOJNENOfNzyDBt+HfvHpiTVNQ6w7k51+i8NJIWVSyyL9rWjpENb+u/4
q/mYMUE+wCKORm5oHeZ7yKAO2RffS3sO9Y+L04RmJ+peYbmT+ZiPSJ8t9KNPRNqdYfwJq0HK+u43
+iRqFsK/UzHhJEnRxX/WOzG/H+qR94BsgbXUNIB9fvDmTF7NPTCdioXcbnfwcrq/Xdto7w9NtbyR
o67UiyvVh132FRHRIWSA47TXm1C4wjwTGKNYeug/QjZsCe1+/s/p6kzXZ/NmTixsbwKABnYi3Z7d
tMLROkQoYDjkMnn7hWvmmdLtD6xtJvwaPGCjKlP1zhbnYLBwSzvhKy9g1tCkzi+6OBAMDW/T545j
KjIasFy42P4MVN7ANd/IsE5WMEXybDv6t7DtfR8vJUUG4fpQzPRw39djPoG7UakyXPPFVbIeL0oW
psS7DdSi/M5mP22Qj1FZ5/S3Z7ThfeNeVoVgxiKUds8O36m7K03USdLHmp9fkU9u4ROjvO7VCP8J
RNHU1GaguT9BosFtUs8Do2KNk6B3SMvHY/Co0GLFu+2NKMzwVgNoFtVe0NVTr40eIlWOYuuueag9
nY5TdElWOvNv9llpcCnYRSHXVFU5vtV1CBKRcuzF4+hj+PtkcX3d8dGnzcPJQNQCePCbtXvFpx3w
oAELgfpqBS5EzsuKrIJ9mMYIj0FF1tXUslp17zoufsKE1sZpcQziFNrF5Ct1wjHq96P2jA42VQyO
7Tq6d2EsCvG38mxblu+NEWAwvA+RcKS/jrsn+8c1DP7syf83nE1IUz6lCxjVQNvn1UybIZyTxUj2
TpJPjZL+9MZMSBckKO120bDZ8hlNlsqvVmuKKwnOEQ/bttRsxp80sp+Jzstg/TmuVXkCBKPU9CRm
6qkCD3RhBXBFdV5SSJi4IdD/N/B2bkjUS6lrdYhKCnQ72TacNDASAyd+1J4dBro0r0Nm+ElQJjXl
96ANg/E1vcRgK2VM78w1We4xSAYtPCYDpHtvhRcednJ2AukNH8RJ35ZW6adYWvtaD9GvPlacN21V
HkOU0O7U4wdCleLrzFlzM4Kl6bz6lpcHWS+xh8QvJ7xe/kD9oKhHqxD3JO96iu1ecPlOHK87UvHl
UNx/p3MYnqn3Lfg7fiNTItoXs3OTtTp8pQMbC3ggod+TI0M1gNDxHjDXfIAnfbAwyZBNkikvv+Cz
NULmNvri3WGPhlUbg2joMjk7DumTkEpXIt8GyDmniccHO7osPF37wv6mdDG/XBmuFWHm6K/Gtng0
gUf+a/gpwiFLepKg6T8XCnTnzMnuCSKO86OCS06j1elxTHFyXvYpQGWRZbsueRCX6kAdwseBTAbu
sOW3lfk8dbmlE8dO5aLlpFsUWvq9Vg6VaznXu/UpP4oZ5eiK9WQ6E7YLFzTQiT1csnZO2HTYpyVA
GCXJBub8wXyS/IiRvOejl/cXp2Z7Wao8EM30Odd51TgEbdUWaCLjIH5X5LGootjGE8VowzCF0Wdq
G8P6GGAUfi8NHHnAxxykNJv78Dqsg2H7IoFPN64K43/hLxb/NwY8IQtP3aRE7jaVAQIYJIK/E3hD
KxvfgDoOALY9FEUDOH0iQIElmKKWseCtS9Uc3UNJ9smRe7GsskMjZ5U9K352aXw2J2ITbWh/mxnF
M+jzFib6BgpIghP0wm1rnO0asYYOOt/aGlFCwNdl/tIMRHxnzN5UbuzLWQYcyPflabq1xiaUQC2P
qUo42MR42YRVKI6o3jp5WhbpK9DVahM4K4jzuuwPN7QT0hJT839DD9Yh0hd0644F57dOVT+lQdFF
2hGkUQV9IMWrGlHfg2KEt9TxuvhGbRyhAtdrBqmHjggmiJZUOo95o2Gbgt1g+c3AEKF7JQ7ONiUn
ilFqITXilvpftx3UdaLxOhbBX9fah5RW7B5VvaamYESyGtBiA+tRi4yufnOLa7Fxwmyj768FLWnU
JrbJ1CX3qzuNaXIwN3C/y4ICTJHFpJ28riNa6VijNwZyzqQ5TlpVS2xkwWoC0/0wOLUUtfOMMZVz
gKKEiWAR4GIGzS6nGowmnk3xmbiR3CeTtgJ/n/zLfZeitbzXmrfUhEWmHuGyh+y+fciKs8xd65Wn
EJWa2avDSoW8eeXn+zuEHJwazuSYGz99h3XwSixGiIBL4a+I655vuRIlnKCpwxVvMMzCo6eTIkT8
wA88T2r5gkYHWziohLYajPMI6CV8/AkKmSkbjKeQnrb7n6TmZDOIPDW5yTqdocXARrZOvR1wbxuh
VNcsJd8x7XnvdAFVWF+PUoziTqC9aJTXuv8dWhssswaEWKY21UToZK3v73KnOMLysNpWDND1zSew
wHaRC/t+DhPU1MDjLDMDCKloGNXesbN+1rP0vQa3PxSxDBkNhBWoUSsoS4yA6rac62ISS/mlwMVB
SRuIv34tcPN09EP/l3mKp5zDC04PhENG30Ro6MybBPSwoaMe6IR2r26jKoV3xeFMeUslsx05QFbB
XSJijsl+ZGDVqSA96bMz5idn0xzJd6EXse/UFKwDSeqD1hyY4pIyPj+9qr0do99ncXDnbKlESFY4
A7I6xSOLob6thR8VjGnFRkNrvf++R0gxAscVdqUuPbAGz5otlJu8g2PB42M1LWb5gODj1EOstl/q
IMoLyBX+Dbr4zXrVKSLSZIe02Fb3WE4XLOBNx7WYuGjndvXNNiSlgzImcnINA/fhZshiuGJ263X/
MJI0br8cp9+34uR1CDcMcJ49c2ENDtauVevFRPLcC70QGmjcJZY9p67xRU4mNPzkWBYADFvZhsOZ
ImFz31gPAmOOx7Xl3wNlUEynpv9Gn3Y159DXLaOMd8hddQr8gZDCuN/9IU73jvdaBw3W5CZJm6YW
ZOT3powmzhJruSLX5fVEv1GAScO5aXy9j2/B01t2lV1Kyhl12zen5azy9ykjNal/FKcYdx26fmYn
A6Sj/zMUo7X/Vbe9NMT/fvQS6tFnHJ1fuJbriz+O9l47zNCI3Ajbm81UMvMlmEqHu5s//J3+lTVq
FzGT0ctuFyL0c92P6W3Aj+qSwpZGj0KNHDogsY+N2zAbj6dMx/xRDJqc8LfQtcZaXc/PTGLk0y69
skvAPHJYs1t2OE/jQ6L+lfQhn07muwbCCFvy6RoDUwcyn+eJnuqY7rD2H7BIN5xTL660yUi4upP0
iaxX4rcGNnQF13wECuginuZ2So4B2ZjPEJxMa61YS9gsyvqe9qSCDIPeO9D5rRxirjxqjwgUDbtE
BBhRfEGe8uW7SUGBbLpFESAcdPF/gJho+Hsm9qiN7T2lgAlbn045BVoEHRQiFcN5h3kwze+gcInj
fzSrklzj3ZH/MWSjc8v+AoOeVbq222zwE0F6rjabZ85C9QAjKvLZ9sPa3B0iwLz9r58vmgl4Lp9R
fZQEaCK6tIMCcaX2hAsc5pxBREpJOTFoB776lbFomINdBTQNDpwht7V5Uk/H+B1Ts3Uv18PHm9SV
cFJLL+wJ4F6ok+f4NaMLdEQ3irULKpFLTFcuuYIQ9YafuAVarfRnKIa/dG4MFy4IazmexQJYbrAa
xuUpW0RcDjyiClFcd9TNPpg3sLMDEd5Yc5iy0B3in0tn9ch9kSK2K3skRGlt6TS3NgSZWPGnSy2E
lEGDDXQJIDBnTQ/ryOPh/uxAZOeK4IwPsnzQR9xul9UR/n/EGhKoNyM+SvgyBNRqXT7q+1w4ZTwL
RSZsPdDHNuCNRhcC0uEhMMyCn2+uvNEkqOpIQBNUVGSIs5A2GMwMZPk5S9eDtrYf7f4AJAFDSonU
hC0akxpPYNg0DqxOCPNAj9cwHIZAMrg29im1JlA9CUbWS4LlumHRPzE8W80iBGrLIgQrsRphEBbF
vitiJxUVk90u/2yHTUR2E4UB6LdshMb/VJ8MwauEuthClVKhsH8oAvhoUD+UIXcLNpHQdMcA3zMy
K2/rGT+MY/WgTo8513gmhtjT14cMn/0qw+ElheeAJo03J0cgYEGSUS4iiZAWQiELUKMEx1HHN/d+
NP4H1tZaabS9WoaETBgDsaZYp1NApYCK9TEKsWAACQREGkapUDvxbeLBGx6OPBSyRDDr/B8Vc3Lb
JiqrpRSK7k81QOuP7hlH1A28s8q5rZen4sNiJIJymp0K7Ckdf/XemzRI2RKQg6bfxKRw0KTVbJEw
tWiIDF+4NjqYwbUaeola4zbpbOEF7grdbfWVMVVM/mr/ikeoOgiy9TJHJSIo4DjYBcns9r3GPMvR
BNj9GQApr1p+xboKRqk+n6CaYEEgEXtFnnvhNxLYhm6mVUfLQ4H51M31zFJZPfK3eo+nzRspEl1a
IQD27ZkLtHEXoCxgaWSNKQqNegHVhSqi4r8XkNSN75Ta7sOwiYEg0vWKX98xQBTQjG1oGxXYITVh
hMNgejq1+rXp27ZyT1Ar5NJ9Bjx5ISZTVWp4/SaiU+74yo+sbZGtE4GIdvP/gNTT7IDvGq/jT/jB
un4C6toN4fhPpkNFl3ezXPp07MCd6Pm1orn/ZaM8BO5aa3w4HGZPpVULaijsGgovxbZGwJrVtgqD
r+L9SR3ocnhmSn2FSVw0hio0ahvgIbZ1F06wdnIiRO42uFqYV7OEOj2qSeBSe3d95yFmcfqFnxdg
TN9/Rssjwa/BTn86/XeIY/OLUnY/nekCb25R5dNUR/CCMZhxwie+3IwAsEckyx8fZOQT6CRIoFlU
Y563+s9Vp6sLZB4GKS7yQ2d8FibBSwW7xuyZXym30pVT3FiPPAzklCmxy6KncfHd+SKCx/c41ClU
+wJug91iu7bNiMP+mfAwIW71pCRWR09USsZSAA6QnFkkd6/ugnO93/0y5K/bqUXuV8VtGP2K1+eN
NntMunepUUsfLhZ2rH7pOG6io9NESu29qOI1cXcLs1OHjZ82z4N76uV5Mrq9yQNJ6zK/PFOYziqt
5NcusGc8l2tbkVsUl9TAGvIq/kvBAEa8UCoCbS/i8wAxQtsLQtPdBbKi/eik1D/5VGOWpq8dcZEX
IjyUNnUtTK69E67+esy74Z8bIalG14LZed4sl24Lo7B9oUSfNXO/GaSOOfkE/63r9jKQS1T/CiF4
cy+Mya+2+tzS1xRsisg2vwIUH/rzDyckdSJquG9yEiQilWZaQu/07MScO1SFUE0EPcVdbzUkBUpY
Ox74ArUUI1XoVyHTDmH0/4YPNmtR4kflqnkhZZ/iLZJ91zG14f3ia0fd+kZYGeWchd5AC9FWwDvE
LhGZm9CKanMzXrrz9/Zwr0i+dWdgln8gVS+HHhM4Z4+2oeIP5yrg/UXa/yHUCgKgsgtVEnP6zkIa
rT8wh/oKs4CYcQE2X45IGg3A2hK6HDySp50iDVw4Hg7q9XI4NHChilyYE0FqeAgwkUr0XhabPq4S
uUpLEqPPnwuNHhQLqgIH5MxSL0ANrEly2Dlkdgf1XeJSu++6D3uNjTj+foUPL+FV+9K1ZzLFlfv1
bRoj6dXfE41FSF2Dw2JHJAMfmu8F/sjhF/WIw/MUkAIFMfIG2EVfK/79fWJX5wdznVx602wVzmS8
zeM8NYV9sDhZcXG4d6cHbkka7W6iXbHBkvSbkgaqXCOnSTmPQ/ENXJsiTLnGMpuOf2JqkhbO7ZIU
s6PPp8LlE0Gsz61QmYFA+c3IPuwUsJP0XTBk0mFTknFHcNXJq8qDsdfdip0JVkmq+Bb0GZOWIq1X
HHB3SEZcjZ7SP9Va48A6wpQIrx7bqO44ezDeL5SxjKcK+E/W3T7E0dUvCLp/RGEQ0JetZFF+dW/3
Q80Gq4DvybtdLfaGkQJWrUEb/uhm0NecEOSqmpOkazVrCG9OLh0Bm0mOHIAcufbBdQyatp1/GaeF
v/yO1HRFbixw4VUe78zx6mWIev80OpfOAeY88iybM9yQ5g+QtwrnyTVOLi+3qT2vhRv9DlEAbZZV
cBRO+fQ2eAGj7l2mlCaZrOVCRv6qUSAp2u9mLsCkevq0ITTuEEGk0AnIFYps+0O+E3FIf8wJdRps
DtZ02seTaoveFjwuSi8DzaCeMGYEMVvq1BiYnVtok2AcOWSFRFcR6st9ABAU3/20F/PtA6CT0FdH
u6S9Whs+erCZ5ChI1SVR1E/RmowfKZzk9Ds6v365co62EpZo1MP4thA8xjf9M7F5FnEaQ11G9Gkp
5WoXLzT+wj0roYwdyZ+7CKM6o2emBY4wPzMGeF3SZCkLbEmrmfer+tYKo31uSNU1dw1LCR1PxZPR
bTcCiuY1EMKGqnLXdgJ/8ME4hhi5C0IBnXPJ2BXKE5WAeTLd76wi9H+WmX1EF7+mYsYXOkFYS/k1
6ifSBkxM+2DReEUbetMA8o24QVKjgxFlWbvTeO6isxA39pG6LwoLA7fIW0HWlCM5ZIuaYi5nA6li
xGhMXSpppmrM6qHRbMGIEOC0pldoHd8XJYi/JkLS2Mdug2+CHOUebafTtFuw+SF00RvnpgtthXs8
IrIj9lcnpCQChp+Lw1qqtXCyo1JBmrl8tPife2bFBLt+zK2zBU6EDQ48ksrSWdMPJH4YssSoNucu
r8TjrfG9CnHb6dLgKBMU0z6KETR8J5ypMtHJYGTuKqyriopN9vpTQdi/gZiBLjvhz9Y5DX4uAb8Z
Led5E04MJXXr4MMzLduah4GJViZgZZK3ZFLxDYgxI1dJms8Z81aspnhdEgRucbRSp6mb24nRAkzY
xtvSoYKq1V6nJGQrMMaIkGK0qTO0zzKcM0lno1UVfe0+rCZM4rf1Pp3HE0FZYPFLV7VRPWZGLYM2
Q3PSGNFI1gRbyxKf8k/9em1LdponodGWpKcAjzjMrOuuKptkNoY1E6grLZ9nWEHoZsHxoE6SwK43
R6EMO3zwNVJsAzgqAaeU0/HyIm6n/chngcaj4AsLwZHKh3WbH3pYmqo1VdoF3iZTG8kRx+Gnk0mt
GY+5wPtCu744gOo7EA8OhEHOPoMQO4w8K3Uv5rPoO+xpRI8A2QcgAMddR9m8O7Q3V0wTi8JrVQPQ
4s+k3ZDnsAEkiPDhQP+4+1pIlzTliALjtAF+fTmz7svmQfXNZZN4k4SKtGSm56Exmy2sSaq5bNGE
iGNpj6d7jibJHrcT6e4XzfGbqeAR64EQTkAa1Ej/LgJGYVumoq3ShS5vjYrbyEgtvQ2TQQzDA+6h
QkTj47ZyNWyEZjKgWw/dh3861fsfsxeozfrk01I4UcXU86NYAC9YyeqEUjTlw34RsMoqduLqxHEn
QutuAwCZ9/virLUXIU8OJgCwgcTfhEnFgbTsrMrtDZ4Y4DRM/5QNGcpTXUq6BTOAW9BnfVHteEN1
NTEaKTElLAF7C5yjdJMb6DqTKKJ4ej2OGTkrem2tdTsZzAAQb+QJ0Inin982LnrzCJ+KVgOMHk7P
rpKBk5FKSxwYAxI5tPHSz668JkAwOSRkZksfJkSY3YnAShvHikBS0vKkbetXA4Es/KJzeihWHUi5
3RQJFIApPA/sgp63ud0CYEJQ5DM6iw5flaazB7f+NniGbWnbhI/s9znyDc8VvKzOYdk9vYaEhjqA
0KhAuWOL0gcSeOTjAyW7c39PxsNIHSOezNFexpsawjWoyMg4aCUtArpwbe/M+pEguHEpBK0rpoPy
uZjF1pnPcemosAxo90JR0Xm47ehYpCTvEl74BziLN0NBNeuRj2lwDcDA3NdbFKZQAiJK4mIRsjHu
LtHS24n2WLxX3JSIm7UU4+T+4JLzNO2snadBNf/NZjmNTLa07d3xIWsNiLSpi66Nu7cktMtLViRU
hlMCIn85Wxg1oCvSE4oTH5SOKvDQ95GowXgF1Se1eKyjuVgYmLvepO5niDNdDoYHpHmaqnbSaKcV
G+cbjUZXHGPA6ygNa3XjnrnXXT5KomJaNKwb0Bi7rQEnYEepWVL870P02xayTG56zvyjio6zb3f2
MR2AryhVdswFJUxiqFowQnACmWyXWvSfsV92HwcrMx/WYcsLvg+fZddVG5M+7t709Lp7nQKhBVZc
KnlSBKLLxtiWVpDxHIYs+ILyzhXm4SN/L15STWtUNFbotVlYJSBcbjF9lT2HDvO3KSHkxjB+ZBB/
PUuJ23UQJaPY8DEt1fTHcU76/DoTmtcN0hysgpIODaDVLzIj9yYg22V4lLlmyb+UGWHOsW8fWnRC
mnV2azKqT6qDbyWiKa67XT3PC4jp2Lynco1d7aU8zJfoGPp4QXbDn75/2YKbj6jAWJ7/5ASuf9st
Yj1elcn58SHvT9SymU6vhuNxV4mR1yMaN0v7/DpA5PvNhReIwJH9GyDBa9pJtKZalLyY0B9MF79p
yUsC7BfXZ3HtgBbvw5dN0i5XzCmSxn+FTTY+6grA3E0YZixypvWWzp4CzHYiG8nkhKOyeVQFcDzq
FIouBSa6neF1PC1Pmtfqz9j2/41zMcZ316Nh1etWRrJsi6aKSzvJTLv6KNoRPylhmWFuvAPZ63YP
O2tz2Wy6bOFdig1H8bOsInSN+xpDXqCCoRfNXuqCFwMeahFODCry4YYlcA2jsJ/Tfe100Gth6kdq
NqhA2R/ioFXU3KvBkdsXuOb/FrNocp3OpRIpgKgibWTnxOnJwd+0+c1cNaylf/x2i6EC6pEQKn5t
Qd6Yl/VNbzRuoMzPvSWxBo8MfLi9433SvpwBpQOyhyGs8CVbezgyVBkYyFaIKHtrdOIZS50K5Eyq
rn7fW4IxGLDLIuslIAdzv195p+XPmhu2B16hC8uCX4eaGTuVQtbYmJgiFV3zVWXWJTXC6Lfxe3j/
tlt95wPKvFW7c/p7n338sWr3yCixBBRcDxaHqSP+tTrOovajE1p1nnlCk+0iAQbjUC2IRfg76R+i
Q/kQTEdDSLBdZk5n8VlvBE94nP2DoSYXo49J7ZlQr9BMoIttefVaJKnZqyItRXDPMySJ5IqB0Ll1
Gt4rHG5tYXN97gq5vGEwfiqibAiHLNsslF44Gr0n1htdP/zLuLg3U6Uz3s9F3wjpsAsWJYRUfHFF
0QnDPQ5cq8G8DbaRcnAvcaiXCc9Kwch/6VPiTNHgX7i/DWzaw2LWcTCrf/T+dzsQ0rDpzJzN+zPE
QZ3OtslfIoVHKJs0Bt/rSld8vRZ5NpwJwfHNiIhGGpU34TUV/wr8XFv20kMWr6tZK5uIsooD4kBZ
9jioxk7RLfRzY/+IX3CKC0jazjhaU6RExTDeoUYmHvTpOx3yj7qiwZi7aX3n5DAsA4yhnB5XI6qy
sgd2PQ0pQqD7xBTlsuWHtYkeX3ABzSBvJM2BozjdZnA4s1S7M2WLDQFGzDgKszbrAHDor2PrEzjR
XZ5zykkobSbu23sph+mSE1RwSo7SmXSttvEZfbVMMLvRH0JR5RJSgZyTeXN8JRvi3JmPJLqwzAbw
kbQr7ZqPNWlapLEKhNNA7lpfUXpegulIV0xW1NMchuGSDwBNnP9+/unsOtjibZ2C65lWYRVfJif6
/AvyUSYJNn+vGHB0es8Gwa0f8xaVZb76eT+BDR6OCEv1u8U/bgOLrikV8SbyAxZA7rnp+t0N3rQy
w5JnBqpkJbaYV2ZrVl7EOjBFfhE4CuUrNqvFxRmJTLMW0lsVoC8x/RvqQvlYxiKbCGeLxuSfDo+K
4RUPbb6YM8hfAVYGQfCZzKTlHcobNOg2/B8mWe1KnRz9rpe9023LwxUNEA8SPx/9m2eK2dYkegyl
6FAcvy50+V61hdsxGTYHvxeoHhHpxRKocvyW94intGaTVMwLPcXBzLOBG+PPkbGDvaS3tTIrenuY
79TXP4NaBMKmrFMng6Yz5GMgLOcfsFg54yBCd+cOx53ROtOi42Ppz0+xCIkx/QZ5T2nl/PlFrdif
wA19XKvdn7b2mGmW6AI/G2VMX5RPXw8nFdkFMh2E3KSMI63usTLePEqYZrmBISL1HEGQcTA8jTij
HKYbSQT32bUkpTCcJTn9Vw8KAXK1cd0gP8S9mgQXk+msZ6QwGFlOAR3nwyKDcsdfKkWtbS4nLJDD
u0cIIWx34ZctgXvxX8nbHJGyJyIgsM3sQbPEwjuVYNoNq+5hBig0nKyDMHBF5XchfsoiP4H6I6ck
RythND6jh5gqhfP4ymRAxlvPpwkzJ7sLzdY1vouTcjssILiQE29f88ttDLOQC9l0SJOywLkCVYm5
afd+LPrK4c/Jy67ylxLZIWs3PswAOeHCXnKK5nlIEiasfMrOcQFSgcqfLThRHW/lO3ir9DcPv9Zf
H/eOQjWWtU/v/psnrdB7eUB2Wb50HTVfKGy66zMmHsccSZS8zHSpN/YRjnDOQkH4ahwRWmJvgfIx
HueuY3e1egtTH9p1N+iyD4xSP4qbNCHhuN+yf4ohZnxTVjZIk1IXNHdXCnw8p7oVZpZ87dkq1Ap2
2x+VPXlpawec5ZoFvfBLM2eFSTqqrK88q7sKxlUbUfWXsjnHtXGp0RXb9+dSfzSmO2ilZyTqACPO
dcT0FtcNm5WHwUGyk8ox7nFP8avkzHj3+0cwHPEISgcVj4z/WSggV/Qwm2I93ZXjdCQ9rGGKbif2
u7aLFxhWZFvO7i1YJ7QYXePkQmm6mScqe1OhfBobPK1jfWEn7/+fqLwTY1rMQlKRVPoWBNuBnRmb
oZSSWdfNXU4DYIripT51K1HHlhHlWMuZSUFQhzU3t9Z6Hx6m6FUq/+oblYC0uMXmfwBBkBeZgoud
zQusQCju9OgwjXTE9atVnXa04lYX/+2/HVImeJffpSaBoc3wVVYkD1ihD/Qw1cwJ2KUpz0agLcSb
K8cP1kFfvRWLgQbW/nL76XDFTvi2lNngcSN+VWD5Z4w2eKSfEO1Yxa2Z0v5dXakJwPRXl+EgIUUN
hZR9Ikvx9LvjjHvGAXww0LBhnrEQa5gkPMpDF4Rw04swWv10AOn14VsjUzfelmAnvLFFH0WBGcMJ
0f3O1xV7+Iam+676/lYHh68Bwc98/YiWEEn4L8xe8IvV/PgNq05+/vnqijqdaW7Xzl6vjSLE99KO
cgvzmNTQ7Pg7X1Q1ptKAlmFlY3fP3rxMHJMpck5fJhlT0742lNWzl9cjdPqbumm3GFxF7hO3DeGZ
Yvsho8sfW1R4xVMe7ZBhgckyyQlEhI3MU6qzBjubbFSWwfNVw1hYJefOC/VqR0F15ihiOjaVvyaB
nULO/Rhifk3CN6cMoC5J/2Y8vVwNu2Gfb0/fsVDViMr5z5RTP58wfx4kP5mOs97nBmiGtO4DeGWk
XawbuZl3zKQi+gta03qPsWDDTuCMRfsItvsv5vQ39WxJf96RBul9MMdR3GCmSuuAgzs2MQip/8Bs
g1uh8SoFP7DyUEZXH86nGzYgBLKL4B70nEPmU6VTdwDxODU+1sx6wNzJUa13BNsR725F64Hxp9Py
c76WJ5oVL6ahSuPVle8jdtYMY/H3xBQcE+AZatEFpiWshkcZMzK283/q6ldv/E48Ah6PDOClDEXh
RNls7itkiRclrMy1d+wE+dFStda63+HGcFjSEswsm7V+QLSQFPdi04kOeHzbdPVwOwC7QCAFqjeP
2SrlRT/JBsJi5IbO1ngcyd/O9m4Sb3pxFYAqd/SrVS6t/WAYmSpONC4y6n0VlaYovfi1AqeKkQiA
27PTHm1eWI5YlPwJ5gzivzDTkEqRt14Je/yVGFb/IeTxmPgtdwklRwF6CUHsknlBZM0wuBO6WMHn
RWRWzRAa5jv2HWUwH+Rw1couOYzc5S+P/uRUvF8KJwZ1wGKUMPtHT65UPq9mdDsK0wSDrsmfnoVl
r7jjzL4CbyZ4MxPzEOR8yxIriij2XHIiwHtELmzlx7Ibji77yAClA0Duv/2JILV2bXq12ESYbJzK
1JmckdMQuF8tqrHNzYvCKQjYxWym2x3XSXBJkQMxHzFL5d7lv5FXr6ZrcIzniqEP9w95fq9h2t+p
S7funuVyBW/T0E/PiCkiJ/HaTKUDZYARH0mFn34UIlGxoTO3jHEp63olACJBjcu3aGpugIE/3C4y
Nsz8fUBPn3ShbzfrTxOrOj0ch2WPl4B8EsNmauNHqB5PJ1olIeicOD/XR2f4C2f70xyUmGhds6UY
Ret9S+50+tPXURANL27jicboPxBCaELtd1wnRKlGJMEU86Lij4ShFvaCtJQpyy0a+Kfv3+msDCjv
TAMbknUbsSSoIqE8eGU6ihrO5dnJUW60B4SKrwR7M7PWvU9aXWBvG9BGYbU7KkyzEHTZP5B64qMB
foFaSEJJ5EAov7axHmpAg3m5qxHdNNH8969MLJEU8EitkP3SKk6ThFKWzFiGN9ulZn6K+T3CEaVO
XPEv+bf6G8t++KskFe2svZIitPgYKUmm6C9YWlecR7R/Cjys7nRxqdZ4k5HeSvC0WM9eSHtXbc/k
WDG6Mv6WTOvww6aQpRp5P4aOEbB7si21JBFY+XaahQ1Yq1u8AdQQdcH80N0HXRAPcnGdpMgZeUzQ
HOXxdPCyjSakW+UwnxSQwM/hCCytfpNtEfph2L/Lj6smwahefeCj0Jsmksw8zRr7MuwusHd1Hvm/
BjgyjxaBSdSMNWhh07w+D/MJ8MN/UZKoIDLy8XJHJ3oxFJyGdFbSUoeZa3xBCgwxRIQo03UPH4YZ
gRqMo6YMTKLXfjHuldQoNZ1fM8mhtL99eVfkIzMY7jePw5oMD+K5pWbkhBkyxuiZwYnrtlDLe3tZ
Jqxs15heM73R9ZZYkGr+/nf+f9hQYgFkfJXLoT3FltWWfGfzT68zA+Szxe+P2IQ4nfNpgX4YZzDj
c2B1wGfgidGd9UJg1OOWCAcseRxNwdGth9BivaAaQ/8be+8YSQJRdoacSsnZ4aGmVy85Q/qfjW/D
npSyFi6CwCFRY+YOiDUP5T8pytHKslZRrlhU41FFKwycaba+qhOXt9NyxXzaQpik8WnzY5PoPhzj
pAk/Vl4AblF99wARygTX1iGS6JBo6TshzyFMMQUC254Xq4wLoSgHd7zgroGIBV2VFzO1cEwDmrp2
dkvYeHHzo1nSmGenbbjrzXGo8qn74Gxx0BTOD5dQIi8tadmYAEGxmjlHNXom80V7YHERDBbe+Csq
EWQJxccA1TUYMqJtDb59sh1uD5mnVJqyHWfgbaUFIcDWC5tml+k0KERbFpuoyoh73wsbYlo4NOMd
ctpWVAZZdQJMK7AT793n2aeDYxfb20XvOFR7bVoIck6FtCGvOGspuGZ6OX0DdddElhoOyWEw2YCa
I0ntnO01k7umhUrW4AnqUwFdbUKoFzW1uKceP0Y05k0n5xEYfzHqaEuv29Ktbuy3hXdOimrOl7Gu
qQRTgFw817qsH3PmzPtBjMrhV4Wm4hsGeTjGP157c04FEL/eI9pYgoOi7mxsFEOp4Rya100nafut
rlTYY8TmFj7RKPOpAE4orY6yBl/Q5YG5ziwdq3mwZiDyqMK+FoSCKQcPZ6DdZZOC2RiZuyVS+Vwk
zs7V8QZtvU0j9Q3hmbeGVpCJ1JYbSmBJlDsuMMokYfoL46LB0t6Fhfx7in71HK5OUVicAan59aYB
mfbBdTiFDuW2V4zins5Ojf8d7xsUkpSOmRp71Zmc0znMwabG1G86DpWBH7rFjy3xrkdiMPnBxAiU
jWtBWCpGoQamERkVUW2nGeXIkBdFzn6EECeAivF5Cl229P8u/M5Wl54yAFdN4a2yQRJ3dtJud8hI
jhbp3EjRlfCAgHn9nJItSKIBDoE/W7NocuAR5crLxrvv8LnqnCCfHbVnRYtdDZGx1nkxhFqZExlc
N1rQTmS80bfcrbuwZ8CEYBP2Nkt4i3sPv5ckBwzVjHeRW9YA+/M2V+xhrKBcQ0PzOUvyD1H7i76t
hmfrKEX+ZU9HG4UgzCZWjOS4RPivsN9NqavwpQqhgG6q4ejxrjOMfThPn4C+jAB642J4m7fyi6YX
wzcbLbjstb/DG9i+99nFBCuz6KuRtgQNea9fBisJkZTVG46IDK01aBCHh1hR2dTIlROflC2m/vVO
wd6sOuTr1NvXE2AJOWSbx5FEWdsh5QeyrgtYSck5PTFFhzJ888J5QthlGfyUXJFmPHclra5+a/Kt
4rEcFsP2x8G3wyRWDaBOFOu+5k8u3E+CsVN7VqqxiJ/8D5m0FmGIHIbcDQDRHsKrXK/Y7eAdaF4N
RFOTLd44t7ceYsHOmOGmacn/3HLLF9g1PB4ApTgLTzesOdM3drCuKnfcGMH4YMbzVtVnPzbMRRdJ
h+Q1Sew82oRuAophbVFKYZcR9bBV1acS4Klj7L7F5tLb+RONVUosUfnDB4hO2UcYJ5/skdf1/381
u+cHZp1qpM1E+YhilQ32iqwHblqeE25aw3z5o7SM7jFAIuFe+0Vv4g2lHcYBHIEfZNsOAFRDKite
dqlqGmq3BZ1S845lShUs172Yh1Y4X8rcric97iVD/JXO5WpWaUNEheHoqSaS7Cy24lcJh0bVsfiF
aFb9xAy6lfhLFGq3EzTR9lOLcWLB7kXsoopX30oPwln29Y1bHkgCPNQvBtwWyvfYptON76CrNe0V
lLwmgzijY0Jv1gjbSLqIwahWapokGZ10+K6bDLQwZGzafOcGxxedDmJpKwsuMpQ1Yfn3r2edWmrE
h8btH+u/YLPUnjbfQXpM81H3CSOFSrnU/2S3GlWsCRyhe2vjK8ZvqA6PhXPiGMPq0GpPqIcYLJu2
OTgLwRBTKgnYbuMkiues+22DFGnE030C0YV46CRDaJBOfrLw84t8u6383ii9p9h9omjqb5t1BaLN
qGi9Me3yUlbxPj9WAYZaIZsbOv82QX5jvInYZawo0bb7TBpPK3CiggYhCvA9FTCUAWFUwAVpToT9
7yuK/3IYxEUXIaDGY9J6qmyxsl4gwl0p+hhO85iUujWqoiHnJ6crGV7chKFWZVHm2aRfr9jsMTYg
3k5vyhUIVuUZaUmxAEeTFnAKkltdFRLNkns6B05EI8BVVRg0PNr2MlBXu3NloQIS3f8Cd9dIO0BB
owptHWnhT7Xu3IOBZ82NuSx2N9C+o1LZF0Ale5/zrvLF58BIQtyBrRMDx5j9isyrAWaYEs3P55eI
5btRGsxp3T90Qb7Ke24WBqnQLrvzHgXBdxc+UcZlUIwMbOH+qO6yekS1c6O37YRxy4/xjeQjITfb
/+AmGNDlSMoQupP71rYg3DaZnmJ0N4vBmUSUG36oXWmPkYm+VuqHmNPtGJna+7Ed9JC9o9UI8dKL
Ks31LurfCcg8dfKhYydHaLZz35TgQNfiejJUthHDqMUaAVV5gMrDZs9HtU6NwpHzSuQdd76qv86F
VNZtx4kt5BV23mTKqjXXm700/k0q9nlzABjOrJ4nmLCz103UIMCnpa068mQ9MuyA1QPLJVm2RT5F
jug69s/XPrCAIXpwdHBpuVUoU5kx6seaTAR3M/la7XvO/h4gj39+sRkhgXKQWffchd9tL0CA7MCK
VwOmTHRRiwn4kMhQKr1VmPO3xJyD0ks1qFX31PA4M7TX5SFwiZuImyRPxOPQQVEtx9pD7Q75LmJS
lRxBrVr6klU4dB69bFo+7fms1RF/V8JuebybQdalnrWcR7V2XPPVNaDQfhy1a8euECZgGZQijLHt
qdZ+6Pj5J5y/CGSJaEkJuR49lI7JfGbreJpGbLC3vZex6jtRfm/mMJ9x0fM98Subw/eOr6KCwexM
7TgDcmtXSaQ+M+rMzpEHW5NFUpA1xefGGWWZlAdMwTOpWqZGjFryWmWEKZvmf/6Gf3BQYNm78hqw
ekCk5Gsbeed4nQjY6Uk6yzUJ8zlwDQO3YOJ6Z6U41j01BRdPyfmb6RSSDI7tbmDgoZhD7zirP7WF
rAZkb9kQeXJEPVfXORN+lOkABip7cVH4WO/KMvvfQU0ljcXL981vGjmpDQivjS5YHeCC6SKTwP4h
6XqWvWm/juWZbeA6JzxnwAWDzK8gwGDv+dSueCc9VDisHl9Y5aVLbQNOCg5R0POZmtRMbn6YzaXv
sbE7Vs+MOMbrL0UauNfwIZW9nYH3gV4LDxqE6sv6RkMv/ZnxT1a5Sk1xxrp/fMZcEPmRHG52pJBx
NwARm1gtpPJK8iThtnHeK0SzjoBEwoti+UYuZfIOb/MNM9bejhYywUP2aJAdxhY2A0fQ4rIxN/K4
f9hDn9tgx9pgQGzkZzjC2AD0uJpwVqgqt1zyO94HW84mjt71Uk5cqgzDdPDmZY0qDexE5wZ841Da
QgT9kN9cRNQIeh0QvICBQwpzyTco8GOfRKlQsn7Z7m7ee9sBtDTPLPy3fRxpK3eo4OC8TXEPICNi
BZV4IU8yuqRqgfbpyhDZ87cYlRnsJwK14ZgJHNB3t4ankfcICd8mM84gjGCqhUchdeBHCgDnDk45
rFNiulJxEi44PwnG//eKdhEEv8UiJ7XLFm6bL0rIDdIr+rkIn9Vdd7/edoj/sk9FszB3k2ZVEjsv
eaHR+ut8q5taqEEoKoykMJZLlpdY2EDhH5zn2vrc7ZkEbc7XDg0prpHFi9oSuBDbAy7x68l/I/WY
9xyK6GN7YuQwbfi/JQkY5Q4PyhiyZCYoVvbbQuR5FYqoSXQOonKNPuBSpRZjxgEPaVCgXxVJfYYY
7uAbx+yETGE9aJ2NA+S/8HKqvE+v8WjHnFAiz7L/bd7kUoSDHuXgk3SjYh+6s/DTNGK7Y8lopt1p
Bqy6QS0mw288YNYnhhkbKxYXGYgAi0DM1BQAbek1Tf0AIoX6HGJCceWms5P69ocGDb6yfq1jB5EB
nqxKCowazz+M3oa0aXLUaUcuX+73/WbiKxFsVWdHWYqNHzCoI8vASNcBMZ/zue/zLAaOxXYVsS78
WB4HEO1wYkIq3+xdj6Lk353AKeCeEdSUaH4Ige5JBjkatagy3NiiW5psLFInMqRpRUqUG+4BF7gi
QK3U0xtFhmB8fnlkEoeEQTMsZvBuakK1yUitwip/7suiswqa2veZC3ukg+qBvGovg62R4TYV1CK/
UNuzhAOBs228jUZ9FjqEEAB31m4r4VgDisKUIkqVnLECGOnUNMIOR6DexqtcYNTqPXkB8ex4qSXs
7ojpc3fvlVt3/QqgPtFbMIBb/gTWGkPTIwyIt5WVJRiGGtvnITJO74NFfooTcqG2TRWg6mPH2aEp
gC9/+hs+fL3+xu/JcThgmVIQhpvCyBnkjuJXorIAYJj5uoquipxH3jsCS/EVhGhD2xDEymzbuMNc
ZUs8y5iRZmel6qtgfgFVJwetb4IqbkJ78NeWR7xXElX6WJDpgDsaNZ5HwDDMDF5xbuBqfIo+eigr
6ChiB42IZp+fMxH1a6Wnt9dePccgQF7g5vH4f+n0lVF0SqRoOPVGtj5jfLzKkfBtzPvaJUPXwiMV
CKg6JaxhG04fR/p2ubMj+pljGANhtm8xxDu2ORPNzdkSp3oZ4TNlJ8/UqfUkjHSApSPw2P89CtHT
dod5Ds8laOehjnE0a+fOoAZA3kNo2mf/V9t4fD4OnCQvieBCaDM4zo6cb0XVL/wMJkxTbtKRqAZt
kBl3+TzW+7eTXqqWgeJJAURbx4s/YsjPHvg7o/m9UCes3gAc3RWQikurdVPMMRIN7Mjbnp8ENMBQ
dNrUtmCEM6tMOc0dpaQXd8g7Dj3rA/SulsAlbAdPHd+IfNTQK9Fy6LSVwGy98Dn4yEaHXvHs91sS
CfVqe31AK/O4RDuNkya47Qapr7rGYMVhWdLLueWYwlnGVjkdGEYgcfv0S+m91d2wuThdULSDT1Vr
hJ/fY+xflG3wT0Ng0DefB9F2TQ7Lo4QA7VfoSnvrhSN/qRBQh7WpmPah9h3BvAyKhUNNhSR4Guaj
e+MeuyfImaCf884DK/9ZuhNcaHsXcni0q5F/c5aNBAjzTxlK2M2GxNjbb/OWLmUqp9C3yvHbrhLf
XglANbVN3IwjRkjYUridR72ZuBqQDGhdFk4zKKZaXelogu1C73Mzi7VpN1skCiLbPnUA9Ukojyb7
KlQv+z2QI56XJDwdQU6sb/GJxZs4KWpEmlBRvCa/eVKEpRB3TkOpZ77rsYCi3tCQ1bOATsifyJhW
LrWR96LzVzJ4OyDOleahtqZy65zPw4Wbn3Wfo+/qoZIfddcECgPyKznHoU7Imxqho3HQ/gqD4sDc
ZmfTHKCink3XFTESfRccReODQ6PQRFoUgoDDDq9U0M/yTpPal/U7wvos88bUzUAVik1G3XH2w0n1
BRYBawL6OSwaXNASUq1jyvHLcMvk0JK0vvMyW3ayYKYLdmYvkPODXqNlpDKmK4j6GqD0kHkemVCh
sX5f+9vdz/EvbbcTDw6GY9a+KgOYLQAmUeN3AfHVJs1ayuZM3IrMCzv13PjwQ+JTMi9poadMRkXo
7qxPftUICW3r6JZViRJk3xpiHiBEvfkx2lTeQ0RDpL3GTxeu5diSoqcHIEh2v2TyBS1WNdEowIvX
cUK952f+MQmW648CYLeVvLn9HRc8InTMNt1bLqDw7bd3CNV9as3cf2PIyQiefOMpgnXS3IcamFa+
aw8Rxn0u62F8Mxx6nn3Gwx1e5xU+TW1ccpFyximKvCW62aQWjX6zr2a+Ze9Cjb7z5iu/BMbyG0G0
vTXD/ppi24Z2pGuvHy9n/PAoPJnWluXYVYZLcRsuU7/FRjZ9L35UA+qhVLlVnDI5NKU+ysAUz5uP
oDPEpsT/d4eI8kkxP/8rcJvePOWJSJVPXnjwEOjQ+8OsskXKl/nGUQ+X+VtS7aJxr9gNjQFUU2Dt
qzuJblV2dFybjmsKQMTtPA62C3kkIRwb2MQWdT/O+9tEtxqs/A7I80/f9EJCJ2wYLXDyGwJpon+/
sY4nwGvYxrXaE9CoJ6Jm3fLaGmZYaYb/EonrTKTk5/hgAc+0iQdAPIqsj+knRMUMvFqNIxSuP7SH
+dRkW7PlL/48yvMftn5P8IBV4GXd3UNemtJtlq47aEj+aJhva5JneHp/149QDGQodnOlUlyTPoF1
eiiQZ4aNIlAu0eR9q5ZXXWwED5gLGsu6jYNMrCE0t7lmZ3NuSai4PqPKLEYtDG7wg7Y24cE73SU/
ewpnu5A8XMoWMiEywJq0iWYwRr3FqVljMQf4dRIdqffRg45l+brF6gqXdMFgySBM66zDcsMfmUub
lZ8qZZfE5SXgqec/x8+dYFesXg++gbR42Gwp81faiBmvWyRwn0hHR4LhyxXa6UUzz6xOak2xaw3x
vbba3oY5kXSE2UTXr6WRNgh/IezQ9SRmvmWCCtilMgNhfOGOVNJMOO7zXQTZFKpy6qMsN24Ww86i
X680+nYjJs/9GLqDrCSj1QMbN/ofZWtoRxFh7ZSyqrhocpUTwGwDomDVuyjM6Lm2EyvDPUtVIBpy
x11D5N5+sUTY8It31hppBEi/EWKy8uHyWq6ZWYtxD/R56q0074uE+Kf0p9IgrFhiLKCwUZQg8vig
hxdlBWb2MjUUQcjscFdTn0P60396EXJGZzCHxiqzJJf0OyPtjxv2iDDCZk5VwxciBkyOnD6EITt1
jTwibJDJ0FtRPAJwGZQ3OIk/6O8f6f34ctHoCQzV3b4wt0Eu/bvWrql3Pp/Tj5es13lolLoENeYM
WUHNiCWT5ja+SSG14s9fN/td+KZzQvuTacu5lvNlh6rd4jNqQt1lYNv63zZwFrDM6kWnMWurh4wA
Ycc3+0A6q2XTGFGxT+Ek7BSLqBAYT0zy1ntZ0q+erzJcP4QfCCWGzYp6QuwJEtsm88tHNjipZzSM
35Th515k1/7lR5MNGoD8W06ONdGtbFKdb8jtP0FN9vHy0OX7+JsiQXSr9mJJasYIjecTUZ0Xl5EC
SLnAb12e7+IBFzB4/oZ96FYMgPgnQlLf16ztLTGD0fYRSHGdZbEGFE8TDS4b9t6liPt0F4QUxPG7
4yvgK8L5rWFx3rVLrJ8DNXdggPxwsJ6q6nTvhhiecYzfNbt9k+fR9Nx30DpX7k013BhoeD9rMbNL
00/0hDuVEg91dY7Qf2k+41aO/jXN98YPuIA4cQUHwcVn0ToQEQBwrmW43vpBxf2TSwtVYko1IZfc
28ApmNdl6FEJWczkgJtru7FzSGFho/xpwdOavkqro+b+wiii+HMLbYhZx5e3hSQoLWcoFLD4jJmE
pTHcxTcI1OStOHqzItcf8jh6k70VqvkGhZbUy4IHAVSlRrLzjFSNQw5mh6Gz5996vnp7cOveGMPu
goJJOrGcgW6Gbsd1944SkQBIOWeoGghxOVM9j3zIUIe1S3/M3HL6XlxGvA0aihoxdkNd9xj5q8GQ
pWU9DHTl+0yG3yzh0x+KPQ/nK9/SA0j9lg2+8VKOB18J8Zpt80abQ9AbLg/EdxU01f7cWiNyq+ts
P89FvnqxIzIC5S0aE3KYTrJdJAM1ErxQsGqALsABwTA+oMGDHf9fmrOt01VRIUiZ4L4LG0L0LfJw
MEKMxsbdQJcy2nbm0kLFti+iYowZc2erEdZlYVv+IM/V0a1LUgvBkaDkGhrx3JQHOC+7FB8V2uqC
uDCpw3frXDJaR7/EqNQxdajezfdVmjhK9YM4q+L/T583FrMqhPrPf49oEzCrlG1AC5fUjy39MG8A
H7YaDKaGwFLPl/TCRZD5ry/UNVac8+NJNfMRQRZJXapTvyUYV3eCLlLQINjJs6oX4kiW04qvmSTQ
xeGoo0Wl9eE9utybEUznIW5/agbqQ8yH+haFEP6XcpIb05p/vwCky2ePJY2u+uo3ycXFTcnB28hW
AtSGyni4CU9VWsvRZg5P9e5ALVWXxdIIVircUfrcIsv3M4Bj6zLVoON6g2drr69nY4WlDUqo5mSA
IdnoiGWLDxTVZd4QdFAEGohcQLE5lg1AGgUqch66YI03XnK9+B2WLhHQCwxC28P+MVWpYjAQ3ZVu
GiRdsDcFsASnMvxjqCdxWJwSmqDzBrS2t/H/2A0KzzYv1DHu13Eee6KVSZNJCgeSRKSpldf42XVB
CnNmUQgTDPnbeDBpnOLJnZZ0Rk44xJ7sp4XiTaG7DRxDodZma1f5nNP95vBCwovRhZXkpw/6o8nu
0q20rBsyln6geB1KzRhD1wItJp1yyq77dtu/uCR1bSJkLHG24ZnW3azj/SNvqIAbX00P7DoAOAlu
k41GP8f1NfGNZj/0jiKsHQ8BCH0WI8kwZOB+7TJzgzOkUvra41cGRxtP28IwmEvYiQLzWr7u99Ex
Dd7i+mJCljoun3yjhzbAybqnn84yd51lnVqwaQ0QQxVlcS2nGU12mrDnzbV6BF3CT9AfMJLI+pMS
M438cRxJOc6y3IH14EZ929wQa6VRAKPMm2HKd5GKUHk9xgwdzcS02FURajKZysAoEkHyLX7EUCF9
7Gb8j4gQeBDQw3xK7O1lB4ghTUBR7Fz7V/BdTpo5SNDz0ZHZ8TV3ihiov/DsPZJzfHM1Lb2cjtJC
0lH6kjs9CH627mnAe0CL2l7GgA42VOxMC1Zc2auFHbsUOgQ7Y+399JZAlutHBQOnXCStxiXpYrQL
m7KW9HEl4SsjnlGgbhvnu7ZCD/cWGF4fvujprGbt+TD0otqByxbgTvUCkVGdwo1F/u5InRCjT4pG
kvIRhXRvLZB68Pe/YIdHMX0tkAs78vmMS+v1EPzhtuDMfbnOsMhRW2gO95lYSU1cReGqJ/ZhOQpr
ZfyeQ+LdxhTdB1OL/Fm10JIQQy1L+OqMbnXoDD54O3yzGwpuZKh0A1y8nm+pGCMffX6BHgIG7lyP
i5ZTKs+uBf07ihXWvZP4+aEaDLeGw+69s9TJBHpsHFkSL4peU0/cR9fS3FTxfnUUfd0BVy9drBY5
NlrnX6DSfRZrxqGj7ZnYcoAs7pY6OSiaVg/TEqmL0PV20FTyXJLRY3+xlPyGgbqYNawy88mmQiDB
Xoj5i6V10MztMnNtSBzkrQ8UDPCMoDtoMf8nY9oWaxOBcBMyhqvyRc24ejYpTtnubWlumFyxyZtd
zSuGyfnedcaqbn8ISDJL+iRSje6ZFOedPzQC4vxFtOUclJlEfYHgWAsYr51/xilt1qtDiMSvQZS2
UBJQrgaSxnk9NsKqdMiFRauVPL97MtsdCNE+n176BpopNyZhV78gSk82111NOl93uf6jLvLS7d5W
qd8Chd3eghtR70IALw230rLfanq2I+QSHCQGJoVM53j5NOJn4yOCVphq5C2PEBvuVNyz6C3Jii9Q
pRQnEIR8C52SVS8+3r9wp3rxfMW9FNfEYy2fXE8xPCBgDHJ/4WF+g6/4eP8frTsSQWBlUo13XHH+
nX8ne+sHV8mGZqNFgxv6ermjXJ8LyOEB0h0cprj8yz9FRkcBOJw6BIlQnf/DABb7ACcpkk5LdrAJ
emd3fIMGaGhW3by3eXztBKKCtVgfK1+zpoXr6/6frTWpFjLfenGijbfV2ULbkJX6rBsHNtIlOZYw
HS2JTj+EOn9yIyPCwhBUAGsXTz7KEnkOWNb/9fKVnI6TDs1PPkqE0MGzJcMRM8S5DF+jPpCNVd5O
8Ch4uK71IPhbL1NZfBxIwSf2/TpXopCkxf56T9YLNwbQaW7GDO9SJbefR9WTz54RFp+RMT+3tqUK
R90i5ZqZHm+hepK4knR+ON1AdK/9pJbjDiQXEOInZv/G+IVXxHrG/VwzIfRRsUaZL/G+uXSmBd2P
HfYc33Nu8fDzsp4k7baUJexZ88RncP3ao0CcCBfdTfVnf6JBcwJSKdNOsXA9LiLpKc6U9MS6OwO3
Mpw/VwYxmeqOfQeR6RngNS/yCn8htmteDvqhDhWD9un+IGkQzKWkxaB3F5U8fY4qVxdGK/7qZw8p
SPrQbkXujtwTDmRLopYDpUbTqJEV7uWyFwN91jNidJcuCL7KTdJKPpMsRPUSFjYyBCSXv9D1eyHH
NyNl3bPEfgxb4oG0GJWmK/4EMonYHsJmTk+1RRyhIkFkXqDeDlwFB3pv47rvsRRKMBB0lUbiE/Fm
q5NPK0ZUfyOzaJbVM3xJGEud6H2cHWU/9c/5dH9hSsOLrWfuV4hVHq5QmKBtx8xRd/aM6tAfQc9Z
hF4vB0YUrho9w1dpmMcZCXsOX8jKrYACjmjBgx5lJW9cLnogXjNbZFs62rS8+lC6jYKQoH06+Ij/
djfmbKi6x+8YLN8dF4uP27TZeQcCL9MN3KH8iYntKWEspdvTBGij0Ak3d7hRxbCV9qSMr6g9SpxB
kD/rbIIYDsO1WF7M5eLsZ9Thr32bFNikWk6V1oiG/0iYK+b5MCMz4Wh3r1d34xfNlXzxe705GjEP
TwGLfqfEkMPCLazh8n2L3I758e+td1WCJ88+FlEXTs41rZnTF5Xfsvxh1sxMhEd498uN8LQJVz0D
6xvitrUBdFN7L+pC01MRAlEdemLXAoNmFB+fZPu9LSqN649b4LXv67WHrI+3xf/5oDmXREqGpniG
u0Y3Rn+jRl89KARASQjdF8+ukhkqS82Sf4lLmmw4spsjGw3a+KxhZhz4JlKCZAOUnbrLUxpm+S8U
335tdssVdsCUXUO0YJ6zkOQaJ6w0iW8q81u/IDfWizo1uptaUnS/VTz0hP9ziI3igaRZ01PJvf/R
Ba/KFT0mHEe+ESwrlhetqBqUKjmwls0XJ+b5SziKwrAmbrabPTzaLdfKQz5NkQzq4fp82WiwLMVO
tiYHONBEcWeVZXMPp68rNteoXuE6ZBUeSSQC/IF74kPe8u3b6o7UQVeJnybV0j9IE/vpKH0M9m3W
EaloRp/8wNnCfMltEF2aITOuA2BZdrjWgDtYqiBR1/5k87DkpN7ED+r0ZRmaObqldWoNH+/7QCaH
sdDEk2w1YYrDvddnKUbR1aZB0tnRGBXHc4hqlus7Xc6jx6QLbkvm4PvYZYVNUz+ptn+2Ef3Z5bEU
74TZw1xR/dl9q8/aR2gGGx8iFWpINWqv1p/TkSN9mh4vR+/O5T7qHD8qCCtseez5o2l/205ScW/c
TchiHD8VA9aWFdBi22fM2NG1QrYG+dJPCAly3URahNtXmzEHK88jdX6g3ki4VcdL5OV4Kg0H27CE
TgM2Ughe8dmidIs8/wCgWwCTcyEBBACR0zfV/Ih5RdEqcveLZ9rEi3AVqGlKgOMTensAxmYo5JAX
99WgPp19iSQ2BhtZV5vjjtfEfstbb2YckoFR4msIM8QnpiP3U2KAZlopXaxM+FEyLI2iwKbNAL8A
dhS+Ua1V4jBrkgQ0rzqUHW3rLmUtBkMuACZ2bFWTAmb/O6I/7MhggcslIUBmxFyFwsRggCNl1Jak
ZZGIrtuLjtLMVLbf/cYZi+0n37DARuUKEY8gdwbASKXLyJDUjvYyxA+qH+zvc81k7SS+DVfQsYOd
aSMfF96/zJtoX3KgmdMJ4GFA6CsFAXoeeTl3803NlsHuVzu4/91yp0pb6Q1SplUC7uawA676mSwq
LcQB1+CDJvQ4+r8DJgc4H5OUNuhyZc3bnnlzXgdVwilWhCmvMEvgGZ9hSgxNu16AG2rwIc3YDcOw
hwjZ6a3XfokR+EYEIyp3V50qUyU12MYU0BZzZHFKi6CcFZT2BFvSxOnHHRfYc/GD5DijCrTpSYN6
5MTPVUzNEaUxZ34VluU3RqEcAH3fx48Gk9uQHmjwcxNBqJIF9i15n6hxrQu+YevgxNWtLgKJqx1A
DJa8D95YeZXGs7YjoowXzOWSIof1nLn1I5M7Agu8/mQZ97cVHfwR2/gDGsDVoWgs0+Xzga8u6hT5
oznLI/yz/ozNJ1B5UBt6LzO5aCejulIOF9n/dv1qtveBdeA516VODEd1Ek6QgxAjEJXjbTvcFZFl
ygkte7IgOwckKAOLXbSpgfkIna8reFHgp+h6X4rh7xVHbxyXyED0h2KzzGZqE6VfLr980NgMZ/gw
SONjORixYXnVIDm596vebh3xDmrVK/gsqfPzzNW+gDUgAA3s3eryZ6i5fFvReXiiCiER7qbH7P+f
h8gYLDErkIZ3igPYMgZm1EmfN07GVfRd7360GMF3uph5pIEYDa3y+LPBx3vKkErdOlAFWqGkcoSb
1SLgSLtU4L8FL9p20RT2lD6rcad+8awpRtm/rGOV31qJ5fN1/QC3ExKndoaRE3tSTfMV2cNcOZsm
Te+62VXvqovODmBFFSrP6CZ0offqrVU5mJMaRcQw2z2oKlXLwD9lE+GBJM6nmLO3FPwePR+JtCsh
1iDrLzHAAUbN/VYV5iXBGS/7olmy1NHXkqwNV/ONY3eHs1nxrCEWN7o1xHM/xwXF/we5KyEvMCow
UIpHggP3AO0KuJUNBbd+9uqBMR+P+oLJPxp1hcAm/Cn7ZqSnuZ+NyQE7Ott7/vjkH5HaxOtcVv3A
DgITsEHIE894Q4KTrZekgoM9zdov7gNHE5A0S+4oPLFuAUQ1fYUzQj5VKEoIxmbzMXf0TALAERKK
3+qLh9QgfakLTlM4J6Tf6L1Ob4WS9BTt8g6QCy3iRqk1zvylOe0uXgrrNh3gMhPufgtwD8RRAeVS
K+AGf8T75fRI9B9N83r1yFp9lkc7DmQ0a6/KDKqo84dyFhHl4/76i8U70O0yGZ08FdmlmeDcTfSV
ZfFcP3sDJx4YyDxw1SRNNorGR0ByYMW4FooSitvvQihz5Yh0Nve+IfW/kTHn/ktv03hZN1jMSmwj
6BQeF/9JdOLfqT5eBzF9hLs7qG93ZpgX0qhlHNh7MRLGTXY3exUSGeAckMqdI3LS91YKQ8yK75qz
6Rz/Wy+h9zLG7D9hEkNfH2YjAheduPsfH176pJ07ypFGAJb8D8Q/xZASts9HG2Jh1l5w6CrD/MQE
TlmFMH973B5gfGR/CVUspx9or0mBzxfj+R0WKvlJNb79b7Bp5ehq0YmYZHlrq0Kc8KGpB8ZfZI6M
VOUZw+P/DZc+tAj3gwg6TMZdjBeSWEGq8MxnErfRDqf3Z5RelOOfn98w8xO0DLwKfxcwvZnw1i0t
PnAHa4lLGHD26votFEg+ozj04jE6j4gehcgRsBIxtqfP/bhIrgx3UycHk60+06jJ1ZcDKhGkq/TI
5rv+TmF8We+89cZzjc+TYlgnGpS+k5UoQpIibEyX9/k0QJG70CLOaLNanAoGjVQkXhuEmps/MV3n
f2zE2epj8f20Dkgz41OsWdyVUODWQPbOFc4vEaeqYInNX8l42JKw6XxWcOYrMrdvtQ3dBUqPRREG
SsQp1ho/EE8r/WN1v4qT+NSXntR8/NOkVIz6EGGup/pt1t/Kqr/6ZysG+HK0HMiydJuDUMhcvcLZ
SmaKxlQ6iqDCCuDCPwgqydSQIdH3dn76UNujjrHOfs4F7dDaUzjWT+WALMdhkiSDsf11hIb0fwLZ
xKthrBxns526NlghMem1JEajois8b5fZ29sFIkipI2FjdGopxb2YUJwxvE2/cZ+2igw+leJEd5vI
Q5Ru+24Es2rmz4vSa2kohgbgdgneHicqh2aql1EdDgrKEXW2NE0jvxn9fIaRpM2E01Le4C4Oywg5
x9hcpewxjYc/DJSYMIDbREaR2H9/uzymqmxP5CeUsps+Ez9y3+zjWgVPEp+TtJWDvaze122Pgzh8
yjoi70OBXfDmYvXv3eHM0BWXapqyUhsuWuVqsfAHukNPqyFIgAeA6hQZ+t4cpv2+0adoaMaYJCh0
qSOfu308umKsFqylbpCQNONQb/o6KWoN4ix4Lm19CUrL0/zYpuOZkOpX9zd6pwnwwpbJCfcfafck
O60C6kmnSQm8crWLlDOGGgShtJ3CJEz7/tXQhznEkPKvy2vdLpX/EY+2CiaD5Y5WxFS5ABMSYCEi
Uh0fvPwOcTrGyJCuTCF48H9B4OMorGGfAGAiHH9vOufK1MOW039SLbDB9p8iCiGLSk3IVBXHuski
7HSDG8HlV+QeNM2fMGXpDoyViGiJS+hQKBr70akhB1MRqWA2lpJPfUITXti0ZfxRdPKgV9DQ1LUk
Pajfu0IRLMYlXQhjUcvSCsthqTgTwqONapV6LF5u813IXbIQV2cg3kW93X8x4WD2YVdX/+6Tx0mJ
Cen5Yt3Vs1tn/X0/0Q0uAggwPm3AYLBfExPIw02+Li5GIUaxm3IOlFbzE185E0GbC9/KYHsHL1Ag
mCzk1NiDaeDGq37XzdVnVBOjqh0zB6JUi1Ol2LeIVS1BVnKDWsSQv0UUt8auev6Kh75Qt0kiuzPY
KEXN9MSyPz7PvDFFQCQfYOek9cvrTntPgePdXU3YLwamyg/kpEtDaBG9KH9UioEYGbsPXLq6fufp
xghcf85wgORS0vwJp7chrqhbdIdoPFH/H5TuX9wVD4Lz34xuT5F8cLkem3oqxDkD8XMHHvH5mP/M
+pN5FamYSZpzP7dg6f0c7ZbgH/zhmc6nPmNhhECLnxiVHEWHoVegrzd6Np8GcNZJHv/r3Ie2vpeP
E2vFB+Og+tLUXAT34YwDVQ8swJSyV1Ka7biz0Gan4BuAtybXAEblPOnOe6yYJVHy9tPwgykhqOyF
4xfDVuYXggmmns5QNAqTi4Bm3svW5LkYnetFkAsIicPziojbrPAdKZ6oaXTmxywZEPUOljGMs8t8
oYhd0/zTh/LO+B0gnoV8CctA9OBcfP5BK9v9X+KNj1kvFHQ94ZrVlu2DNugmV3CiaQ4Q64Arq21f
dbb5KU6CZInuWjTy2eTZ0PuLA6JVT5mpZ40q2Vgi8+/AZqK9FJesl5yH7WteGErbPsh1gbcnf0Pc
ubj5ETJr7+gA5UBYMZXCl5dGiWDobXQ/83Cc3bg7dPzVmxaxO1PNE2vqrok/62gkUiplGgiW59we
tCabsOWdljlHGULhzRvf00ZiUzDGeLUdeIaKSCTZ+OcEjXYwXMuv+A3HR+2pnlnbLjVyuEyzMuVJ
FzRrvKuV6ArLOckd6s69BbqJ4dezRZoxViHHpReItCoJFKoxOxb5F1VXFgr3EEOozanEDl2jyJdG
8MkOHB8FAu4KPzzjV6aYcfBybL+ze537L10jolfLmqrAglxcTuU7qeey4g3HlF1K1MszB+lShmRQ
DL0RXLQ2FtGIA4tHqnU7/zPDsp+Cr7XkSfQ6dWi3XPlTB6XokeJAjN4K48cqZ2aHhbKulNmsH6td
//2Vp0gHFclke3nimEvo221qo9S/hKU/gblc6hTqNMdmD5T6oTJk0XLUuLuFJ9ETAet5RktHNWwU
zEB5vW9OdweQRZanItl2d45gCS924oD36X6O+Mk+v38vwb4ghMeMr8Iun32cO98XI3PNS574eHcj
Y5tz/MRd4QbIFSeG0m9lhWcmk+twym7QbI3fhrKA988+AZ5SuNYa0p25ssUp4VNrm6Fkj1Zw8p+L
/S5VF23g1cU3jY3I513RqunM6VNuez+PEKK079mcnNVmHhn1KIyPAoENqRKl99JQ58VR9fV0PCi8
Y17jfV8Le127iE8BFxwUKFUvG1OoZRmmSsWXK3MTLK8RsyjNezD/Xp2zhGyLlnE4pTMejEWJwSY1
Ahl5lvlIA83VapEPwU7OFKb35zqE56v6mVc32xfpr2KL5qZ51SPp53w4RnhtHxFWx+px32Y0dNki
qR29pAt4YYnoDWnBk5EmCLeVQ34aPTNlCNSUv49WVx303uOIWM8GF6b2LdiR90zLXl9S9gZ/rFzU
pwUvKNcNvnwQLGw+qOItqWCFMZRf4RVwHGTLSKQD1g1NJMciuWJz5QoexugyxcEU/0pyYGE0tQwz
qaXDEdqKMIhKaxknZrdHdxJuQ9Cji1FN8l4bSOo2Cq9C3+TiHMXMfe/+kkHeqdRO3kFHvk/tLgA/
d+flRnMkkE+MdF0uDPv/J+RJ/xybt+Qj03IBQU0XNnONdEp4zXhTivi07oPfAuI2Rsbz8GlH76TG
ku7BwiwvYaNhxWDbYou22sNFsL/4hhY5/P16C8mq0c9wDJ3Fi96+PIkFqL6iPS/Vpb5Kv/Pek+Hw
PLgkRIJwk3F+cXYZR8WDnHX3NPkijwCj1zJTlPLvuz6WR1lgKHD5vDBEUzRRm0IE0i4PS2TfGGa3
mf4Fp+hH6vBhzH4Lo3F73w7R2c6D+7YP2jD8WySOmN6Un1GjcbVmF8JjByQPfpjvGlbXYjTrAxjE
4zw7ceznOBvaqQYL1oFCteykkju1L/2qkEtqbSa1NY03S+xeZ9a6jFB3yZtyrJ6Vq+S+tX7KgQfh
vNDpalO3a8KteQn2uH7y7gat6SDUUQK5uPRhC2ff21zsAVlvVs6gVViIdviOFucnRDZeAtbDomof
RKvH6DLZ4wLiM6vM/tKJaBb7+ncTzBpBmZ728SslW+KfSFMT7EJH8bK9PIHx5BnjWHw6OwZ8B6a/
kpYAXE6r1g7dQYKZMjQyo7tnn77OPGFuMiFWl9auAsOl8YBZfDn4Jfd86qYsVym34Of11PgprL5X
ni0alhWJqrjfriA1wz2U45ZBTzORLDrYF9kbLD/g2Cxk0EIWBeclZgxNvmmWWRlJeTGUUHJl+sH7
uru2On/0YAbmRQgLijAZ4ti4Wgdk2SWLoMZUW0+fHvxPFKAgC/1jOwc5LI80V+6zaOT2/zX7pkcE
Krc7rRZaq3IJjX1nqdYTa9QZYX73jSm73OETLIn40c6NXRRVyKrmbsN0HSgxj0ydBCjJxhD2rZXX
RHfZxP2fhqPZ2j0aDvP0ikpsbwPJh5PgJ7wipkmUIRA3xsrpRXyayIJh4wwzX9uw79uFbgeCptPO
jGqyBKrHlRNfbngecPmWN46jd4V2+c352KliJh90d6d81k6bI+6K3LnSDGFgaAYKiM2Tpg+WL0Ya
iW77IkaHsNQ7NtclTk02pW5RFZQxp3SmRk6dkG2BsS+CXL2KG4CTnaBvhwATuOd/TOocOSetryMm
UZ+xRsYQbIasEo/WnMKMjzy63yiNcrssXW6KJC5I/L7eMtp2isE72re4DKLTKvvD7kZy/YaC3Xum
rmICmwn4fAV0VcRbj/tuE5LMS5gJ8MStZtcSCmq8BpgFEm40wfaYsR7Au0xctj4Uycr3a4fkEM2R
8usgJ7i8Khw43AnJh2f7Fz5p7DUjO8SOyyqgFWvggTRj3h/zAEps6hNtXvFuaQjLjmiRYetBCBFH
QA91WGncZp2hJ7on1IlEoifSnvO0yGVJDEzEhWJRCJPB2ZKHIB6kP9IkYeIF0QoumrYdXe+KzfPc
LSws4WFGEe2tRL/ytFcN2/KQ6qT7CT2uu8aNyqE//kpSSlAeFZN0rqV721FnpB6JKh0y4aIDgtxK
G50CY9ePg766ZWz5TPIOGdWEtsLK7cVEy/n+WXI8BoxVUDf72G7Sc3b5Al2iZRvAlGhvTwt0/xqr
xXQRTWsv45/mAM/nN6ohmiqWDh/rdEK72+bf4UArCmO9ON6ukvdwQXCdEOrJvrgLWOr6Z3Ga2GC+
C0gWbpF0cg32ZINI/bJ7ltMa50VAO5AJjWGFeey3wMmgjnAmW2wXxDBiFm1O0CW+ZD3pK8jJng5C
+VIBzq8NK4x6dg4dhejQX+lI78El4q2TtX2ZXC+APKvZq6UfVvvUUR/G6A+sO539VCz1PZBAKjCX
GytR1en8R5ir9ZF12qBK3+RcjD9Iz7JGkOcTp8FMuQTUwlcwBq32dO6Te+SKxs6PqZMebtZRm3MG
cG1J6Pu1DhxpHh+HKnBhXiUCSFoQKv4K6JzWgX/Tdq22XnbuZLfpMMeg8RDa7DqMrBlX7cG/C92s
V339RavpaZoS0fw7B7HWmJ81raeOKFckcWCupZvMVwznnUYy4EP/voBqca5x1PKhqCwgMk3MrJZI
ynEvi5KXcxbx7ZrfyYzI2QXEGaswm6Ffx6ygkStjtHQgh7zyJehgarSCwe3c/MLp+j9Vr1Y6C27G
XbQ2WpkcaL06A1Lpj07rIOdDJjZCFPBGdC83e1iJX2gQ3sAR1FgN8RvnDmQY1pYkpxjI1aJY0cHY
/mSSOZWHNNpfn602R1n2ZEbyZBRktCeoydEeqfPwSYjy/dWSD5I32paluDqBhB5XKp2dAEFreJu0
27y7xBBVPUh4ivZXucg3EQfK6uKzCXpluCcLfzX8HI/rx32ISAtsPU+LVOSwpmu4Ah/PEncnH+XU
TwpX90haPhaWeAQo65PKOBOvBXkAYNcnhPQ7Xo6dTwr3O23k0WDPUzqcVRp4pioQ9xA+wn2mcthi
MWq1sx78NY/G5S8DwQXlpsczIngTrMUznNY+4g5tFUZSw4d+RmeC7cdBbgIT7eL8ZeqMx+TP15jE
DtHAnLn1jcfgTxg1Os5CayyaGJdJvR8mikK7eCz/KVTCGSO8OabfgfUrVKWSgZKSI5Bp8aQ1WDZq
h3mq8ovYwwMBBw0VglnzIm8kZ7mHdcc55uToFuNohHNhPS1oVbX4DfZzQvYP12okax5M7lyYuc8a
VDf35/NNnQ09pVt37qPuxXGRLe3IrRCSz3lS0SH6GstvJ2e60ZTTdZcfApegamYoSbo0uyX0kPqF
QbVPQq8gc+Ors0i0bOf1rIoiVkdWb5ntfwlniWOv8GuLNkOq5KGqlR7SyFzOA2oyuj41B5xUoeZc
zN2RefUUF2Wjy/8O6hsisLulCwpRkqhtHsHKGJ5FFHH4HklfzrnJqKvU1R8XIAv/+i/R5efBLM2u
IxYWjqmdVkoPJf2K9EixCW0+SoN89KgdKNQId0GqaOzX9cQufV68tkPJZAZACwexlGqYpjoGx9qT
s0hRVI0+MxcFroFdGvXb8aCzUbcNQzgy8hw8cPGDpmUMosnElelclUE3O2X4RP87WTUu/GoKh5UE
qT5fIf1HATcVz3jhqap+f/W68R2o6iBACaZemQXbuaEKfK8f1D0v29Qcr09c/DUfbB0znP/lMsGR
bFeYxId82HhEJMHeaGb/dtFpoE1wEV50g790zS3cF5toGN6FZXhyPs2TNtsAyEU/idMLcgmFDC/J
RF8J7bs/cM73/vYraWY0e8DUghe4gzRDt37JpGOyFZgb3pDIYE/68dIYpJgD02wo9+kcNiOz3Hd/
xOweDCSDPHmqrYbO5tbpU093QDMREs4sHG03tQZ09idmhStE1VT610bDicreMf5ilbh1tRfYUkl4
OVjkF+o35tRjQbl+zIp0HEpmZO9Bu+/aATGBUDURojPVYJF4OViLin1AXKOJbpWd0rDvz7FSQgUC
feOxuQOatRk3ZRhThoNjbVkpiTljrzxTT1Dh/CMJ5357clut3DkLc4fvfPleis3ARh38z/0YyUtI
QVLtdhPy1QbJ2pt4L19KdHW4uMNBFxN/HL8TO9SOfrw+67FnEyLvM7QfVuW+8CoScrXmsMMAk4rS
KuF+jjIA4tnOamiJG+DesysOolsgrbEynimnY4PcFQ9jFz8bIBEwHL1N+6J9SGFI2um3ufqqCO/d
ibARfjw49ZdxC+QAWQvIg9QfS+1z9B3TMkLc9tErsP1JFj6WLR6GPZoDwyRy5QfwLciOxs1uuGPo
e/TP8SiH51Va7LSZt2r3/OZE1NOXIdAZjxlcgyCvDTfTNbT87BRyJkYUD85MmtBETBOxUNQc5UHI
gFliq9e+YBVbc+54XX8GIS4TFyfw2G1Tmgq+5A9tyAglBXdtmDr9Wyn2qhxzBpMXUEIkB8Dz2wj2
u4iSDJzEqPgiMkmq8yt3BBdGzSnk29H1MEp/AXYMsvKx/zDuCtP5EDBj0Myg26VKhDwT1PvUxs8p
7NKvYm0eedsCkwYg3A9yaElka3SZs9HX1OcxuvffQ3dfshhKIOJSd8OrXKk76lyAfJGBd6qx+XKQ
lXvpzXiLggTiN1gkECfHuVUWE2Qxogvt6YoKcraj5e12VQrUgrY/pYbKayxsivmBKdKxr84iQulU
m1toFfWuKuFC3qwuQcvWFDkcEqFTiph5ePeOH1Adwo8DE3vr73avrxvowKKMbQRlUMXt/btUB+7d
GhG59plW2HbteDCB5zCMC7HRbngPcAXZiRHZBpXbFDftE9AsgR5Z+d93rpsxaiXdJwDwUUwY0g4N
+0nGLM7fW8zzZ9+lRYsnXXS2ukpNDFHDiKiFZnnT0UqzCZi+rYSqIubybv6rgVn6G8EO1d+WWh4k
qWieK9+0L0d6VWPd+oI3gVfI1+s2JhjmTY+3bNeLYGeQP49SvW3IaDVn65csG6lSK93Mo5oCmtXK
xl9pDo6Ylx/B+WtahA6R8yeMxuOO1H7xpKKkISwD4I2+xiF+de1Q1QdLboWe8tcY7MZ76LIfJo7B
UKF4PycOt7/DX3cMAiJ4+5GjzKrHaNYhYZAj06ziWPczAR1YHX5rnxhs5PJ8gN3M6XTYWVLjGjM4
W8gQwSv6aq4AA96SRnMmxcCgQLumzoxH1rnylSLESyuAFNv62+r5Y2J/ryw+VOIoXF7chbDGSqoT
vwg8zIGathE36vsOug/wJGUk2F/vuZJp/gEPWa+Ux+5PtY64AoD0ZW9UDnEyi1gn0u7DUb3fY2ny
LBvxW5iPRUYpxY8QywmSG8/MxL02ufJJa6Avwc0MCmBRg2FP1n3AiHYIik8TiQmcu7+XP8qpXFZd
FC99/T8zW4ug2G68AwRacefvj0I6POWCoHo7Lqk0ZWbyA39S1LHKHaA9p8B3zBXF4zL0ojTlqWvv
dQzILingLWeVf774dgdnb/cxgn7qxlENfcO4HB2OqrQTAMFD4ELikWAle5hMyfoV/NzKjPj+MY6N
DqtP3l23JPomJxEt1hFBhHcyiin45Q47t5HdnkEuD9RFdL1/FOgug7ccOG/azvO/+hAdfUndSaEa
a+DW6X4b0Ks+kqZZLKWg7QaepXJBM0Vboo+hIfDp6Ko+5InnFu83jZALMlmqdQDdgvJUZvn2AmbH
i1CO+f0XQmceZwUP8b3NVB2rcmnltqZj5Om8EUZLum3iGA5us9Ryxrw/mUuuxfC+DrD5pbPFI7tL
D+x0LoQ00zevd34MjFMzxJeudNGKUoZdmqGN3wIXMsbE9Nm/sOXJUJ8weDi+D/XBLNAduSi6dGM2
wbtLHdLnuhDD5Fg2ypv9tk2LePOv0Rj73n8F7+OtZ0ID3urlxi3Vb0KCX64NGXijfP6D0DLrhMCB
fRR362Vr2n4+VZjs+rjzO1fX4kdTDowHP6o66G5h8kD91lmIudUIC7b99nj8rMxe6A0PtwnJJlB8
j/OZ1J29d3k8qSggegGak4OTPRfOLuEZzhOV9QvRkUbzWalOveGKSz1f15vldbUUNv+CGmOolcG1
V4WYFvMhbpydb/I8gklxJbSr0Fm38ArGH0stLI75XP7mWoX/OOQobLrVIm+Kf9BeesFIObLRikHV
bZgsOnHoSCJFlPdP/SBYfpUPBXyxOYQyBwnzvtvsS7VUsXJs6TBHpq+ncJMhIOx6lfx8WZesxHCi
LVtx6h0SIUquflg6T63Az2LYJ7jKsqs+7U1N62wdhPmXr5nhbNUs0XG3VVv01Tgs5EwGvT0HlAo4
E22vkE9JxXaVinpJPx7pi94WiVuwSdy8x+ECNhBrv/KNerJD2KI+GuZEZd1DsdvDZqbM0UOHOxlo
UTmpnEMeXyYOroy+6L2VoM7uCnY72O9vYObOX9Lz1ojxnMugYuCLzX+4EKZiQLiARqZsNpCCi/vH
AqGKF/X1pte3fQS62E11X12PFkKMe35O8wmlCsoMWU2X5Mn/vheDXSX79Ax6DK8LMJ4prj+/0vlf
nkM3ojEvZAEqmUtEAL6+zvg1/NpYnvPfkyOSWsmEYIH0wFhvCuzDVGVPX3+wk5yuxcUtaU6ZWYPa
T1yhtBzHFaEstSTklpsNa9vA7ozwRcbZF1w4nPfVKpVEF1QgIpYgS4Yp1ZbOU0LtYgJkkLNuvGNW
Aa72shPfQCdLPnHhcNMsD6VBYHIAgFFpOzCuf+hfgF3GKsoXZVZOQiTuEkEYxlIFyY1sEehZm9P/
ldc9GotdBDn2LWQqZI9T4rXK1z6hHQG7ccm7GWLTqAluXAbqQJB+UJfuTwBSgSsmt5xc4YRbK5B9
KUNRXnWPKJT7bMexwtWtB0F9m/rc27Naaye9tC3h0CbHa4OsKHxSJTUcZgKZw0flo/HwjgZrVZN1
jg3VGnkX8VAodOKQ4KtnXA6AwNb1T1uHWbwEhmvKw4ezHYP5pqbWl9jHzJdIz4sCZfYaDLLfdieD
jgZqq80w6eCM6wQv2FALLQSqLJoDyyPKE5knFG6dLp74W6VMUqvbCZ+oPJVnvS/ahCdz4BAJebEK
WrtOXybjEVVGP68o8VwIj2nIoduiaBu1zrfamV9HaLSkkTzVrWoyZModh+c0wRycSTxzowW2nF47
sczQcFKCQGH0vw6eNsGYORER5nDB3BALRE255DVxu1/tiGJgCYMHCvb7nXVJGmSrT95SKjNxu5cc
DnwtkSKjZyWJa2rZ1MhA05HH7q2IboB2komptF/mq04c2bAhAo2dhVzpcEV7YNWG2oxUR89WR74b
bskeBZQN3hMzGSJWS9zflWhPHbcnd5Sa9MXt+H0ibB4m+PX06xW1a9iffC+q/O2k7BgmCzksqFPV
G3pqcoQImhHBQ1xc5P8IjkcTNSIfziufPEM5/10arQULmDkyS7GOAKvEsCMOmYljfugWc6VJtA2T
jGovKybVPPaXX/QpI4Tv5mmqkUra/Dfgr2RFboJjUJC9CFx0SbH7zpJtTS8pKX+8m9dp4XzhRXYt
Faq7I/sngQccCPX4Vs6Vr1c/xlY0fVDTn4lTzXx8FtQw36bRSawYclhgDZO9M2/boDoU8+MxWn6o
AtL6E/YIxl5d59UMXs75H2AcJDjrI4vELETM0EQCFmOVJ0iluuHc6SfpJAd4/hKA3g1fWFPG0UnQ
5XRp/dMQkigqgh/GyULLu0ojXS7oUL9IdAxFNqcR5hSQ6RFYJP22HXBW65fCSzAak2r41Ys2oBEa
g+71lbnB2eU5igppSB52Tw1GrJ5MChltpXLdEXZEK3LpWl5GnJXporiyeAUBaprzVvo9TxWxNnEE
RJr1h3gu3PUNSZX3n6YurvNJYwJAe4R9UzfA5j974W8bW8nvGhSqNZYGu8oJ9hI6fdCeEGeT6i+m
GTz7tmm+JjBWMt6QUnO/OeYjHshOcE5oNaIpg6A5UW7EFlOsthz0MihSecSniU0kzAwYqde00FKN
02thsFqIwpl5kUHpEPWIN9ldQu3I813J/qHpd49ZzliWgQfDLV3m3Kd600RCVFu9CgrtfV7vR18g
+F462dcuOOKVu0ZmiKJHcX2Hw7zZDw1sKIiMVzIl9vvUd1I/CrBCrVph9ouIovTO31/lPP7kIkGN
psXEVcmXla7MbLEea2ezAzafGmqqxBUh0esiuvJxZv+kxNgmoR02i8Sg9C97myW89zhpfMmMHKZy
CEE7CN310zG8CyzBOrt59F6iiRhs1RRUJ1pTbtHX5dE/IZ2lpkBi6flpqZoiX73vH8qTDQE5bpiZ
gIwAznXbGFbb+gO4+5Dfu7evxJsny8AUNoa7myWelbk6wUixstGfrFG27dlt5IcscFqlt70Geaxe
n1Zp0RxZ55L5rN4VViYneiZUuJU0uWX0ZcDp1PvrfibC69wPEc1zzkt4mlfFeHxmn3L+zZNvSjhJ
bQYSO79QhDUt1SiU7dy73XJYm47Lp2eYDdw6Vmh/FqzQdx/QlY17LIG5epH1WZj3JUYlIKuiXWsT
sbHUhCPfw/gU30F1UEZGwdoclBGlI44hAlVyA7+4SlKFxyGLNqnWLSpSLJTJAqJf7cQcmtPmTZFv
wqy916sawKxi4WJ8YRx/AlJ8F37k7sIz/vtTmOb/svd+EH7+QTJA8zsgQLGuxKRkKwkD+ULY+sLZ
aPlz5UBXnoieQxMfbMJZXCSN0Z1ZCq9+wCDke7Ho6NZPvBjkLAHHYqj48sxkm6SGev+I96Lr5mSj
ErKidRops/TaMGzAtjU7689cLuKimMpa4lHmqpTGXCAV2MjoVH5CNP9OJ24VpN9wfApb+pymTc2u
RGnVREfAgND4cCRj61xsxEzye10++KbcGxXXtV2h03imvt76p2zE4tROqSe1o7/b848MUZdB3sP4
wrnefOFIzSy0UGYQg43TPVO6Gak4x/rTVJnkhQLw6pSRwqzx1wllMVKja99erONt9qvqcVrMzc+C
+8MJQcqnHI+45AL/dk0ReSvuw8Y615rfWSxbhRnLWkJ1XxZOTz3AIQfOPqImn26GTYoPamChn4Nw
F7VbKozYtubNuuDipdE8CUIaCxtMz8GYQpgKuLisFbza9lGYSrEFVPWJpmjR6AtcbfRaRtRsWiau
Xgw1VrXxH0b27KelhxYtGl1njndxelEDR1tQebEawh9xz2h70CVV1iKUkGe3DjA8kdO2BIuHpFNU
4Fe6ZJNF1CkRGvgkQoyJote4dwnznEm7tCrQf/AhAUdkeimISci4t5wfYkbgn99i3mpDFP6t43Kf
EufvCnjse64MWLzNC2Tm6NxoWRaTDrR7EXVdYhh4IVtbunTDEXcBwZ/pDrM4rwR8mbckN5/MtVLd
nTufgembfRn9j65a2xqT7b9iYQFA1SnGq9AGp6dRVCT8psLvjl9Ve/HJWfHMLnIAqGcEdTuxcsKk
1ZS3PgmXrr176nnDQuWkjB7QyXtFv4dlxLTRoyqc0p+wvGqdF0e0SCZ+Mh0Y9LHjAvPwcud4P8jW
eHEly9DDbiKd95Oj6XcKfGt6YaO0BK9+kbG0bsgBlt84eZk6plHaj52q2zY91ifMK+7v42uFe+Xs
qlabhCACJRlAkqFhygKOBLxFT50VK6/GJ8MMcScmkLNIMe1N6JmbRCpRncV4IFtAylTil9YNjZiC
b/SZ6JYB4HssrJnahUeXdjBcfqt7YfkUBmsRS75Ez21hP8nxfZhNZUg3jPgaBXl2PaJUtyvLtyEa
9QL557yrhqEg6v5hZagkboG4zJOC7YKMUTuxrqLMXyC83osgN9S/mqSym2IqKnjIbw6dUljPClqW
OtkTznQJImmhVFOOGH7FcwJQXRvIzi0CPvpJeKZ3rK412/vpG2YWeQ35qwWLiJfciBs7WAZKvYe2
6YXPxCoGiKKcqFJhgRvCMsM3g/745Rn0XowGhC58LH3s+XjjYgW40B+cMd/IqaPpaQe9SvzyLicc
KYmB2ByyV0iWCKJiCMJ84ZbVUiB52VRjD4JRXUrboWpOV5wNby6ma/ruHm8WdIDEJ8esESEYlRCg
MhVRpLsonCKh/oI+rtYxL08/ira3Pi6tZWqsNrJj+S240CiTvQ54l9z4mV74cV+a8eU25dufTxWT
zKZOY2ovMVfG8Hl6yDJxTCFj21mJQUu8+VdGXMg/a8k0DT8M1ufXlQDPNQsadWQ99sOdjhi++6nX
PYErMJF7aNpmYVXszeW+/IsZJ1NCz0NVRBG9/9+MB2JLhdXiu58Fty+1GVHXJcJ228o9tTEYs7Wn
VUJMgBN+jU3On3+DRJ+dZcmFCBIIgi0k8AQGpuTcKeJyE6vaCN5skWn4Lygo0HtlzhustEWMDgAp
3AQdRD0KNNgJHJ9PQvVBT3RuD/ziGFKN0nMqUWPcs/o9SZfIOEp7Xk/vbgzUi5VDeEbCWYHooJcZ
Y6oInzdvNa9aBXWZND51zdi7/S85dbM0++MfCYeTiRY3LH9D+GbqkB/WW7Yoj2MfyYFqcD8Ljs5j
wiq6WUeSX1DDAycbHUL+DZ9SxdykfWik6kHXy1wFIUr5jV5S6ksYWOL37CVoY9grFoJa+bSdA6r2
dUFomYrr+etKDtvLVOQq0uNLnm/TGA1NwJS0+rpQf6VvIjZaByvguP6lnEoJ0YFjXO30qHB5I/aY
kLBIkMwruaJ5rYpWUxUDfycRKQ1kdNXt2+pUAVbPEE8breilpOryh2hqJWpMdpRwi0+VDANf4VYT
fDKb1B22awiAl2yxuQVbEFPF6oEMkPNxk3gWPbmICQFFt2B1qq9dreIZNLwjwJScOUtBOPHfnzA8
Ilnd4pO0SiFoXxFIULaS/2B84vOFrYLZsqTt2BhSo2vf79A6n9LKXIxmlghTA4GtbgBJU6xvqXlj
YJXb8zc4agfl9YyXdjxWQviXBsyMpGa1/UmEK6UpN2gR7nbLRyZYKGjjfqbonKaMZhgA9uP0GUZA
7Y+tDKN1+h/GA3i1woP3lRhJWGjh+Jb3Dm5VisetxK3i8OCqHv5oATkBLeBljdZJdvSOJI7nZpNI
Of8AYctY8z13dL2rLdIEvwsSejA1UAZYKK8IeQQlgpq/w2cVilQFfUnhVesvWnEmpdCN5aVqmJ30
QzzmtDY9J93WcPho0+/MD7XEYffyC+n8Zdd7I6VamrCnX+ZAGUTjHdeQq5h3EP+FNVB/h4zuNiZN
bUK4/G8fClpckQyJg/IUqfUNdJ0h1fQNUiQ+zqQugvip5kBFdAMAU19sGL/CDQeGb29+gfu36qfO
qOxMqWNzmlCRfZ+YbLg9tmdQ/a9atap3IYnLsPBRVoadsCPtSjSrm4ZVNLOWIvx+4taoSPBnAdk3
5K0ixfm+F/EakboFSAW0zUTDHqfw064z86IW3CKYSnpsZdqr51hr4DJObdP3o2RCGFNn1jwOqQGe
A60CqHpkcCw1EK8Lr6zcJjsx0GDqt2y4Ri9oSHtNmG4ZOvvgApFbB1SY7niECqolyjH+Tc7kJ5H2
zZq+LZZC6PP7RNEIncUwIVsTlrRuEhbhzcwwBOBRd/tIkQQFk2QxSsJ/D4aRWG+ghEgY61KGP4rD
gJDRnxOI/N86VpNxycyrZ6wsDQYcF3trC356/ggJLqP+yulYx1oBCA+K01f7L14i9dNZBDjGkOGU
3HLMqpPFY60AEJRsdE6cqx+FjwSIIM1sW89Ku4+aUFEcgUdISsuXM3xW6FfPKlZKnwuAc6I1O7Lo
xkt1VrNvJx0EgLTBx5ODx4wmn9t2CeD+f4Qt6WvB3FHxSTnoNPcTAkJAm/vtmN+q17aYlNPSBera
CXvGdrU2pWSeosu9HOeply8jrQlQQOprDkBNexhj91VX8Pkif06mg2P8ofqinrzt3xQRtiX1S7c4
1o4eMuNEkqUC6jiS34LtK4X08K99NZk7SRaoczsCAKoKyk7J3+xc8EqWeHBJ86wtDDGaxBKehJGy
uwAooTFgiaVIEuPUU3Zxl5QttuKvg9/cL7ZFF/BUzQnhL2Xg8t+A+GLV14I/n9rfPkvUxCQJ3dLo
m9vTv6ZY9du+f42LvQJa/7W+NmnS78gnbiOk7Ev+6ybyDJpSYE6fS6ByKupfHB6euIPlnghPy69v
INtg2fK2+LVtQ5sS+SdtknQKp3hOEMrIjVMBCoE6CGTeO7cs1bGexyS/TzqnMTVydyF9Ubf5CShL
pSxzM6nxOeLxg9zjUkLgKquUo9Tfm6CYEeCJUgX6XbEyeF3yPv2FfWlYCYWlpcgLqt8DXTtzGNE+
CsPlFIlHzMPV6JUKlfu7bOiAF/2dRJE2T2k8nTETYBeXM/XlmBak7t2FfnJ6ezILnA3hKvDu8XWc
jeDZGEi+RpDde9Ik3TqUpGMAzy9YUiU+bTHGLcX5DNJCzfNkDt29E1Qm6beSXM1LfjIXJlGOrVDS
txeTtV2P4qod/+UrUvnwHWCDYF8ZMz9Cs3F92II14BvB24RDeZExQQ4SCJrLWhWAtU2fQXZeXlZq
aCBg2x+0mX0b4pc7PwW8Fe0FnlEJ6Xt5wOZUbz/uwsFoQMFgjcBaZMgXJTd50MqHvzJfB6j4CGQ1
Q7rcNIyTFbEZyvkKW4Uk3NGxTidE/ut7y4MLn00Sfw27vpZ4OugY7smtXmZLDgyanwDeLEvAn8nM
md1wLbQnE81RViBcDLxewKh6u3cOheMZ9KlomBQGUmAmU+KuL7LOrxynl4Ot1dPWFCdeevYSvM1p
84D2w12wIW27/Pf5Qrw+5OZcV0F0tnoIbx1jy+IPz5bJlcS2Azl3s/jzfnQeo/Ee8K/ss5pAiyf0
sMfbG0SXFEJ/Yy2AuViR5OW7SgRFwi2jiUAP1b9QwU13Li+qLMsiQBGb6zCZtOlLl9gfb6cbI876
lndhei5rwlX2/d7y5mIGwDpMUrC7a3ajOLVKZkUd6YBaVAOXSufSiAZ7BXceLmKV7ZrE61v1naVv
U83YTZa8Rsagttk/6Pk7Z0BJcQWbNl2gNW2hIJhB4FGWp6sVgl50zHbLW1di2IB1GjrfxudGwqLZ
5CJ1/DdjAPT14phx5HTMu2GQzVxxIVbSw8fH7oTriPUN+g1R1Y8l1qi8ytlzlpfbYZKHQTyrCxxC
ijrGKTsajbIzq1rZH1t1FrkP2MATFIRVZGZiQACBy5WYH2JInZYh1GI+fzVwBRORF0NqGAQlmCI3
U0CDtw1e9lPI70yEqZYVhA5R5LeZGUzcd3qET82oDUXMnXXuQiUeKILp5/HnbmC2rrkJQu8vCtQ7
6U+8zUJaoWco8O4UmiheaElH87NSJLLR28mgljKKF0TjSuALRRgMU9LVmAl9a/6NhCf7klu2QUAo
dEYleDdYFq9TL1vSpK4080pkYDxQVKzgE3TO2J1yxYn2vqsMBlsrlfOSUEThxxoVL0wsH2uuUJl0
OBQ+dT6gMjeVfOXquWQJ/w71mQNnz8Eg7JYiyUeg9MJqw3xEykUoRU++/cKt/TKsB+29zi3I05l3
bqtmRZrsej17CIPw6/4pvXFmj9na5TFyYAMVRexDX4TQPnBv0AGqL5wRs15M7dEW+xKy6/rCJUzc
DjV8rJCt18JpER5bNQ29jq5dvxd5HB59FJfHqPIk/Pi45CYR+bzIyFLi2c3MoVQQ84tpDpNMtoxp
0EEgTqMmLYico1l/+EyFM0yksL3ay4r6jW/ZWsoMPTbl38eJrlXinafLrvwjRGY90fMsGoPqkxVl
QGPHfw13g7qYDRUX/YoeopZjpK+ELOOHk6Y4CynbBY9PD/up8AglS7n3R8UAQz8WM02qAD7GV0Go
5ww4N1r2eAnsE07hWJegyquck6rRVHhzZdzZ38yBvePaOwkbKKW/yBzUgEvT6XLO2bNdl/GQEnPE
efEgzrnjjewc8s5Oka/jGwseWt7OGfF/DL9gq3/7H3+GSagx82eUJCyvJ5veLT5Pwd1UMSu49Ceu
XKjEtqgdMU50Kldqk9+VVz2nGSAvleya/G9UnHW17LG54KRM8lT/CGqXO3yIZqxaU2dvJKRYt0P3
MN8qa5OnslBdG5pUnjFYrrt9OvrL7UgfTtqLZ7njbFKY7AWUs8fwylMJhJH5G5TQehud5/NXHB5F
VMxezzeGY//l/LfKPY9F4l9LKO0LoEXEUcoAqEERt29otx3BQhKrrj2DEbQmUL3iL0gNFyfFGcrm
u3qPuwhv2/crerlXc9PEAoA3ZVtqInYjiOkJyZlVQ2QAAChOOio2jszc6rGVsihveb2wNbMt8Nun
PbG5cnVBerv1XXTXPbylVh1X6muFhxq39VtrSlnJ+gdxefyPQFvixzIEmE7zPd1jDkD1bRzxCLtO
/9KAKNQks1dsKUAhNTdhJhQgEVeVf7w8tvcA8GDLFa62ewWP5+nBXe2Daay2RDlvdUeGTPT4sb4g
5wxAstH73ewBFEQtVNeNdorsthjKWApmUeIecw0iy4/E5xQhwr0pe0nFA8+1JsYlQ6JLpaTSwZ2M
qx678knbFqexdEBrqglgcmWgdfH1jYTXPnbdLx4QUYglaFrrY16dDb9PJJ8KgtCs2WHWFEmJKkzw
Kgc8Mzgz1c2CgHP3iyAI9pBXcpaokxk/ivXLAICJucB67WtulHffRNj9rRgKXbkpQdzxIwWshRHH
hZojUkEvA2Tjr417ewF24Sl079+OsVzf099rK5M3twkjcknwgPUzxZ5i9CWdUNnC3SRrnY2+IAO4
OdkAFp7JvW+2FJeaYoOW0IX5rCFlNyY7T43fkp9peO5X7CNvBsgbJNjqRLJNdwFV4H/dl7J7sKxf
Ploen5li3CH8G0u+P6z+U6k1pvZzkiSyaFlroe7QWAyV9P8IR/NxpdBvv4X3KVbvzfSlP+deDjgu
33zheAxsFG/JSWom+FYJacfzPa0Z7JrgOBHqSmxFniw2MZUDeTUJ/PNQzphlxcZ7Ppyj9Udt1hMQ
2Av5mXQ5/iVNjG8soHplaXbyUVTsmWb+ZqBWDhtViS0IXsimHDEThQjmZ9gXEw3nJVgQ3RHdJcXb
kFhj3FOceWHceH12nKQPwhRTq9mNXZ3wEAK1WZoE6c+z4joa7ktQaBO0D9d1WVYvRMCkDuQsqUAq
H7hMImfweOXVSQSbBWc60qZkyFRiuKcOrx3whYq7pt1V3UrLW/ItOkcIOBIddtL2Oxa3Nbvb9l9a
U5zQuZUMYj6bzOmru0/FsIyrfz2CntzvKW41VtXOxleEgCKEPohRqgY6d9mQOqlGKsKKDe30iaw9
uyk97vM72rNTSXOrf3G+y0nwYeWZwV3/Gk/ejp11vU1OrDDI/kh43n/JHgcgyd6SaeJFMg2Vj3UL
l/OVCB3cK/YHrGqQXfmDw/M1vprTvhjR6Pp98WPzmZ44WHMkD3iWzNPwdxRcVEnwWOlIgVubDDIy
Qq7Cean1Rad3xbO2DFgPyP6A88xh4pOACJpDDM4ip0g2R8QbVeFKuSB54UOLufrb3Hnr+uES1H/J
y/ye1nRdHxt3JNU+0Tix07IrV0pldH2yOUrnz55jArnwLd7WGMGBCJEQcC18/uC2qj64JxVrJLFr
QK3U8eDKnAWyL+EAiG1Bdi/nmwX2Fvkd8T0ur4J0AViSSRn07yizd/i/zVqH5C+J5fgy/pE11UU9
1Tlpe7rT4aTp1ADGfSnDpU9QiCXF+iDPv298GY6wxyXd1vX3+cT4cKoYNA0WSGDvL5r4KfLYm/ra
Hl6SHnGgoIEvAorj7c655RiSM8rpd66rhN5Bn6LaXr8CUHdNPugou97p2WBLgY67CfdpUrLGqR5V
2cBP7ZmyeaUVHieJNOMMos7HqkpwSn7NwXC7IiGvWV4ezk4s7oI/dAK2zfStAWz4vn32qzoToPW4
U9ubv1QNhbfqK5xiT9tuhgAtYjUGuqZqtdV5WQw/8WBp4xIYy1revGbXITwDTTC13ecatWuExczx
qCMSBIyqsHCQB0/ZeGEwW10jotezsaJIfKVPqUfae0ASB76yxLpeKRY/QPo/XdLKNC9zM2JMdNl4
mn05Mk12dxo2BOTkpMmX9m6JFAtVmwnrOL3GAnnUhe+2IvAjJ+cAcrd5LyL2wNxKuzwAlluwbl5V
5FletiDPdUFS9jiXK+iuFAqTcwUWvFFNQFAK5W++wr3URmgWQLK6x/gYOrL7zImwbyJjNT1eaRNU
O/Bs2pxnaPbD0/fpOranxVEoIj15ZGA7glUJPV5gxqxs/FviAvuuFgD3o2R2Xgok6HvqOJsPvZ1z
tMcHeuTgStIadOK/Bzmt3ULAKRC1DCpCV8QEzhc4TT+gi2SABPAbcMLmJKg8a67rR2cFI63fGamX
3b2l01Bs8CGAbxRrbA6AFRHZBscU99dPF1CL4BkZ2IgKRs+BdgeffAeX+4ENnzl+kt7805iXSq13
q1KmGTad6V/RFpFrQxlRDWNsZM3kWEfNEmGBFB6xil+2dqnmRjMbazQhJgagfUlfrvTVgI7mPUBu
ByTRFWETqSEzVcRS4UeqNBUJdjcbRYvvfJ/uWwd/PNYDYi2w2dJGHbr5qgpFeQ26+m+x1FZEp1pT
+7/81G0X1IdCSAodmdwU6x2nI+89ar1f9XAZLCKWaUX9PTQ/slttOXOpVSrqnFoCuj0xUNbdFUhh
Eu72jiw+xnR5UCDhlBqaihlIzFY4fMSH36zfgSOAJegpL8FAb4E/gpDNe5PtQ7f8wTbGSL44bFNG
EwIWBrepV7xDZE+n2Nf5aqGDZKyN8DKSzznOInjyYjxD9fwkEtXQ/qw6JX4IidlXqm47hq2prGcq
+J+rhiRLyaNC31RDHE5HF9Jzb3GxTq+0s/F3QAeXLCZ7O0eC4G+A+xmlyEisqwEHHJGx1XAoy9xR
h+LKE8dEJ9clmpWTRONAT4Q4xEutFM+CqDcyeVvHqUkUg/MndMFJAsey5lW4KRpQuXhgeiirJVGA
qGFM4Sl7DlZYC/yRqOhx6GAtSY5jVg7ZbMwvB3436Xm/BRLr1tDkmtoT0jdTeTsrKTRUxjVZDbke
ap1NkfuXZdypDnMTPs9O3JGtTDsrnxOB4KmPpfNZXS5D+q4nnnNojPvBx5Nhb6uY61SMRmpSNMp+
51ZO9rZQ2GVUsPBP9t4Cpanc2Nzesb6V0GUSLWzN6QTwEO2pr3f/QpI0hZDOqFzLqiPPTFHc7nu1
jBiyuO2EwFVG3qXNOWj+jFIQQ+AA/sSc7dbt6tbbzlUROpNe1jgVE5hRrg5VQPH6A9MpgSiYVub3
K/Pe1QgqtvwOby2g9a72JmSfNTbOY9TDHj3W/lsOTLd0Z0eDMpvOFnWgfukkLGB4/iyTAQYY89ds
YPRzarzXIszCBY1rasA4RQao+xsF2Ivh99AhCOCXLj5eWJ3YEqnF+fn2fnUuZkn96HgTJVF8RDP1
VVNOY89GskXv55Jw2+qxlzt7TTTURYARqo3BA99obhkCmOfZmjBAwO1o+lt4P942FgzQbTPeb6qt
IDfo1PmFoclcdZE5aNHC9tM3kZM3PChWvDLtm04M/BgwjbXKESzBOB0Kas+1Ni+fEhtV+SfCmsZ/
hOJNcpm/jLVFQIsF7dpw9INovg2CEaq5gH6hcxbhYqHVXc1sO7fjNgthm5nwnACQVKcvqouJmDPz
UPT/MMjxiuPKGbpd47Ae4hFc5mNJhRAAAlqDB0WdHM4f4q03XpUBEMUsTIDV7UnOvSnSSsBc5u2q
rNnbKz5nxsqwq3bRqzF98/iLRzgFQ3oCfBYYHa5KawtqjOzEbFfrRJbz2Ti4pnExuxnurZEN1tT7
eAwB91b7pFUJ+EqLRhK2VqDj85cPHJo/971Pm2p5sbXo1Z1aIN/WH68zKGMf5DgVY7/tCImjyUJc
UivmVOsqAtV0xEhbtICYLk9iMEohT4HX70orTm1GNZH4i3kcLOMuG8VDmgGPqki2vuoig2Q8k8It
8JD2I0Fv4oZ3bK6xSnrAJfiEcL0yCHIIk1reeFmjL8ZnPby/jElwvxAr3ekLfkkUcgJOcPUxl0oO
Y9wBnUFmiKoRkscFGVYW6KC/tvN/KuZwrRGXakv0Gd1ygvspllo+S304OX/ewGcVO6cJVjhPmCaV
+2K0mfmEbYgNA2WjH/U7TXKiaM4XQXPcfvehFmoVv65/HrlOC5OPBMto71NsSX5rTHMGdl+5CS7e
crUZhJM61JAJkEzXDUMeqrKAFY5+bGmHPahMn+6vo1N/ED85m97N+qI0pJ53/T1RPnNlkDStWBeo
b/yyseCB+fJF+ydzb9MmqSPSg10lcOu7DnzbQSWbYdHsV2ODPhR8QbNCHjOmHGpapAg8WLm0eJjF
Uda8yhy5/5o/QywBwieotz3m/iqHKthn2xU/+xynmGDxzF9vYS+deC3zFeBe41WA/vv9TMVwcIt1
i0Xxu8nTPixYYgZz1Wz76+UrPo/mt1KLmODEZ04FlrLMwjFKAMv+lg754lfiuSkRxcM6S6RRhdF+
Xv9w14frED3uUxqQyosy6RBUy+bdZkqDWmjHBPSrxmMkjYUHzihx9/WQ+X0WIEHKWimnEassD8Ld
fFz+6Bp6HTxUo3hncgXsWBNM+UaBjr4OtuRYSi9+KMAMToDQf71q/kn+YbNVADfYllqcdCCCXzSf
jIhwP/fvnZ3/HoiUqq7ErAZ5blV3JEKb+5Y9Jey5iqsOCUvHYKWI6tL6FvtVQ73gHi8Zt7gK6FVR
5aywjVE6yvKm2+m2mT/bFU4PJ9gfB2z+Oow5R09ZMDv7p5jmcIRF69DNYPrnB5Fjz31tb1vO/I/s
TsQVWeDIbIxEcyk0xFwWmZ5BS2mWFrmQW4Sf33TopFSAwBQCnpS8oBEbfn2fZtURv8RP72oW7jyC
fevgHyF61lECC7b+PWfTmoLZlAcM0g/xPna1C7JY09PBe5V/BRg6bDTmW3u4BCFT4pfCtGf+1LeZ
b7VjRHQIGtetbyTz3Lrum59fsfykIz3YkGWNFQmgUqxPYP/mnvamAs87NDdGXGz1QSomoC4ThdQ+
M9+oLgXQhcO6Mm+cwkRblpFbS8RjR4yLijJb6ophMIAlO2R9I1yNVcFglo6DC9eANS8Ie2wgnUqd
m2RvSYMWT8xQlGhiywiU+Im6Ebj0C+WMAFT9PJ3+pvvLU9viL5fTfRJXn56k5YjzjuW+aLltFzK+
wNIi2Y3jcqWFOSMS2PgHLj3xHaITX8iH/koiMAZuQqjlsoQie9tnmplvuPLFNkFwrPJPmJZUXWPH
D8DHHQMPlQXR4iczYWkdrAhAm3jKjkLMh6y5P0hcZlNPE6MK4G6c/iIWHTH2v6b/w/S8FaNOI5Wh
DDwRl4TggBAKJ+7b5mArtmYx0jhb8s1OSefLHSBLpwf6sUo0sLlK9HXzHJ+37WG4wz7BVH7amTQR
0+zpQV0B1GhrPTBUWBiZa0uA+fzJALwnQg+z4mABiEmMuknqf4384oTBIEF8DaB9xGUaMARdSJ3d
H6WXjpQ0rUHl4lwI6CKJ2L44PVQIF0Y4z6UW7e4FrQR3ughDN4kG6VL8sIFWE4t7LHChFfA+WbHH
VJnKoJq+mn2KfPI+4O5uMxdEsF+NzLMIoOkKHkelceCNsQGNZznsfxFwZiF/Mzvu7hNf3pde06U0
1LXRgIDempMU30L20RaeeP/mffs1JMj01FkMVUl5w43P+ySbNTJLZNyudiIAv9KuzOGLg9I0z47f
WGAU33CZ2kyjdf/U04Kac74aiMF8pOiFdhT8jncnU+YKe7mOUb5DjvFkFL5BPwsdDdRWXhKxNhPQ
cu7ocwQF2Iu0C/q26cqAhfGXASDB+TsCPvbMD2auBGFFpyjxprFEGPdCsYZ65Vc2PN7SPbhg+kRT
WFLMwLdJ30rs76hnwlRV7+T1tayA2QW11/4UDD0ILuxObUkD7IrrJBvokRedqFoOsG25HMtLPt25
t4+Vk15rxbgscijARjlWHsYeMSZzdnYOmPDQMyxbawdPApqCU3Jor5EJUZ3fWD38M8+0Pu/yvnOF
wdezbqIbxhwe8AAUdANjlq7ldbkW5y4gLPX6ulFASShpMEatPXR6x4ZhPYY6FIGdmJD4wBPH87wr
eAHpnO1SsTKPCqiYeKvCelV2mlEL+7Eq+3KqshYGUAkDgo5CBVWvFxvH0cD9M9+pwMyQfKVcmkxS
UvLxgrnFUvx7Vr+xNXfopW8W6r0nM3u4GqEUiWO9dejpdheijEINUVjfrrFW4j8adPvCFSnWMY4V
BRLqCxMja5l+b7azXSWBjrFB2P9ANkQ+ajAGpedA5GLqUKrtYSqSU8LVVuz/u7hkYu/0AOt6ByRE
OM1CBd50tkTTOZ8D+UfXdCjeeie6+OPJgDviLY3Gs4dAZzN4z7iSns0csPGzWEB0weBZnGhI/L8u
RIMxCSgzNEfzwdVvnSilUds9sfeeHdmmlI1uvSDj+tmzPrlWFSQ4oQGcIIoS1D4bDIezWL/Ra2hq
//UzLzH3FlPeA1Gqk93FRy0dAfabW36SmVM36ejh9+PeCSrsmcqFq/gvOMYLUG0WjfvUulAOi+Dh
qw4KrSCIontz8eOzla1ncQnpmzzCwzVOBiGBPdoR5dXi58iZNLlMx7Y2XoxdMQ+wGPVu1ZSinJyF
/8dTHm8kF+2/qU9ysgcUPEQ65yBC3KD5DiX4UUKreNSXlRvLNqWE8e4Ei8QAecAaUpfGOoVJovqt
g6FbN5hpP5eEedIMCTHBnZWphFz8VsMWXBogwsjgRnmtg6SuyDJtsPGDt/oFBPPIUQQI3Mwj6s+1
WnUdz4Ii1F2Wcox83u0vF1FRtq40ess3wNuTxMfJUYfMDMW6TPSfOWayscG/XKs9THIbyNPJN5T6
M9Z/UomyoFTVFeyknIZJabrSRFuH58MmzpDSa4gM2YYGP0UpKWraWnQvNm3QjX7t4uFg4lGJvPzl
JGSNrxoJqAuB8ZxN6/JHU4SOQZ5sQ83fa1RIsCxJVSjb+KN0w3p73CfV9rVhMUw4pfJ+UTUS1/X1
Vzp9dfxTwsR9Mp37ADTUn5l220oEm6rhSjeQsZv4goFgHZr8o/ls27FKXksJf0GDPEmX6mYJ7Y60
fbRPgr5ItNB5j937oV3dIUpuQVDEa8W30wmmsSmh5pNnyJsNimaSyD4amQwXDj/lX9+U1ld90Mti
haRnMTyhXURDnVJELaM7Vq8HC572Qi+6eDnGBZrq/vQq6TvuP5a5QQvvkq7D4WJ/BYMEmL6mz8mA
V85RD99Q1byNN3hT0v68xH3EHl3zINU50NtbjBSw0nuU/gKrOFPAg2R0Vnb3vn7uKlhv6KYEIule
4mlnf+UO6fxiV/rvqlGKCx4mJV96bdSQw/PoeOSKiiyvPsJ+zmP8uL5XyhaRZmosUHnPYa8t1pD9
UYCQQYk5zskfH2ZnvPRNeVuEc74oemUDC2eJVqfzPjMZtNqqS6mtgWdh5ZEIUYtO+/ZjpykIsTEX
QRTFapy50THaVr3PwWUAKhULunCUasVcXVWk07fftinSGLgPvn2dhen0hpEAFe+V+bCuNjmKzDKL
8Jmyp5gQnT2t34aECmdnE9a7C+bfzlfCmr4mgzEyQLOcOLPbwPhUjJkKn0gfy/abQEEG9nohbR8y
0Cnp2P0j5E2WY7VHhotXPOo6IndpNweelGGvZ7Or20xP/R+CVm/QRnFHJJLH2kNbIZqS5Xvh83/u
eCc/ar64TDFOuPDjvVXGjTz+7xP8kxGIpS+yW2u5u5IbwFAUv01L7nXYNuovBF5WQT/KRQXlM/eR
fc/P4nytVM+j9nrIKSprxYep/jVASFnYn21FDSuCo58+b7rd8oVAv4Es4yHIvH00RmOu5aiBcX36
g/EvFDLgBcXsoGpxMF4qqzOUtqwwXXVYRAS3IYiVfg0QnsQOn4GHXMJ6gOyAbGHbCAdOyTq8OIYg
2Q1jyyjqrlb1JAk6DoTTZ78hAzp2kAQH9tc94OhqKT6jzIkn2QRi2KujoD+xnKS1SHH8eqCViybk
736etagVd8vlH2bMDNMngdUoVdq+zhmyzt7iIscYKJBtYEmfJxkZb0n3bibyut86fDMrJwaWVdx4
8CUatJ3y9b8F8twAoBC+VR0UWXvTtMpawA1OSIiGANMTeYZi2yhRWsRiQRL0thJgPp2KCHSDIENU
SdGOLvIQ+K6uQLVX0vjAB+IIm4uMx5Z08C6vOw91nktGtWRH7ieO0qTXKUGBVSpFHzlGTByUAhk/
R/gaV8N8/kDs1/mlUQDrzFnJmvjNu4ckInevGVu/qA4jzmjah84BqOG037LCvs9UeGtq1nAtIJxR
WpSASlqZyHX07JixkjmG7t3LEz0EJGYeFyWDmW8NBgePj4ZM5UxQjIvIaYkSdPVdXzcDuidUKII1
3eFs0mzmf7RMi5gsu4qNJ3pb2l74PvsOQh8WiPpUe+llhLTMph7FHFhE8ArnvuOyTWX+1yuk2vWR
xo1VySZcc8bQ6O1bUiGBPyKuyJXLqKzXjEv0lryUN9auawy/7fFN9wSjFJyT9hEBj3ymsTmXSIFM
MLNwH/0VIamHt9EhTeyK/Qql0/ZD0DycINW3meYHDHjqnsDm+EFmHyUbTNKJ90XdFot8GMPxVjKV
7qumO7Z2TlNaoAVeLb6kJabqgG0qhGXjpTd6bW4ARKt4+RJRWpJZZcRGQztPP77PdjNTB52BwloP
mY16e5U819nipB0TSmn1O4efA7P/CF8ijiTPdk5kM0oiWnCJ8vSMzQfpncmvA4d4GmIP0z3KtnGj
JwqeplipjZ3RdtshfqM1JAiiR/clnUyIttLKpUWomEbNolSH9OQR7JMoR9XjcxcXyBiAdG3Z8xfx
UcI7rRyTyZVRcehdAkGLymdOCbTLlaLaJW5APN4l+1UAd6bhJa4qyPpMcS2ZHf+ARoSkVPwIkci9
08se8IgGYwtRxTGzcv0w/KpJIr5OJtXmPxnRs1Z8SmuOjyW66ZYp64bjsz30iXE+wXpi86Obn7W0
RncpIUxViddTKwXUsBBAw/LQn15PIafZj4fLkHYZcvQGR/Su9MgsxF/B6PpupnIQAnvhFhrw/x2S
HbrzdnACHWbi1Nb/QXYAV1aj0lv5TtESr1uOoZcJLJ3p9yejI2ROuClhaJ8VK/0a40fJPCF3j2HB
YMRDEFahsxXOaU+3TR0juZkXRsJ6raPpWbxWxBX9KFtFSKCEr57ZqFZDU5lByYeOJL5m4zksadKL
7YDVS1sUjjONDseFG8kg6QP23fPpj71SQUyv5MLyKou/5Z1X9oa9cDVEHAQmE9lH3HYYDZDX+vFt
5qgi9jgxXAdPKgu3/dlisiPzKHxsV3MjM5sJ/GzwlUx+oRi61CuUucL8ygAJnNIjZj1iy4omBfkt
CZw1B5ybXsUZNyCNXFlP/I3/T2tPkjX20gQUNyNwWa9cj53DghKh4GZ33xGiJXmJACwwTTcY58ZX
0ew9lhfyXOCNe+INRfcBTsJ4+XB8bxYVrmv0Je60xPEpJha2ihJrhuDe1IaN4kFrIzUJO+OLOq/q
3x8woxh2ahhyuSszEKsCWpF6MCfXhxoGWtHtT7Mi6Ngyy+xX8j3xjF6AHuqRPwBAyxUIpUvGSZqZ
bVvjw70s5r3PPMUg2nsAgCm+fD40M8j7G0XDB5Zqt6ok5rpBikJtAxvSvs4U1l9c3US2AZWrRWbl
/gHrnEhjQCoTxiE1yZ5xSAbWv+lCZgHadDMdrIyAe+nZcffSVIL/yYK3BgKsW0ZQW0Vm8o7hQEAg
NDE8eqaI7TzXOPB6RCb0cA5TRlkMD+DsKnfScZ/ulSfPmRNBXd/UiBdktEIjoDE4zWSIWiVWuUXa
JjZEMtVvTNXtjROCFktsgm9CsawQYZV1ZryhMQEJzb4LgquOTUF20gbZE9VviUWJmGNK0jlo3Ssh
iRVdfY7Nday7/MK7I6O8FK4rmlK0pAV3pfYhP8M5xfDpurg6ZK1ZkiFtQ2HIp081bul6ne/ANRRY
AqTigTC05SROP3a2fyZaY1cySKVxIc+I/EiYqj8JyFITt/b0UpxQgyFiQnEefaBZcAgI3iKBLn3c
BRxWb5FQ5qmd5fF0bqAxKN6+MzY2Wz7eqwDds67u2NZCSvmrhp2noJzciDTS6xBVmdSIoHsmcbV1
1XxpC8v7Cqy0czEdRXQqbLJWulopbcV0EnBsdobCEArYxq3aJqngcVtd5F7SvueUkHo841Z6SUQI
3E26kbTPFYCEuywIDZa5F+byB3k7oQAzkfQdm6agdnjQrat4AR2835WZMWr4sbsc8A9peVFzttUH
wmwYuh+hQaAsxfmubo/K3uRfVbNotuX23n6xIHKCQyC/rBqxKOtBOFg2v8Ym66U1M78CGNJREkvL
zLJ/LuD10Vfxmwsd/NP/esirOFftsn4IPB/QRjBckxOGNMZdRZ2hbfDCU0t5H/xLSywU4HEGCdVj
ezBbxoFhcS/yFMaXfvq/VccF9n2Hh0tiJmpWC/M22bag5K+vrWlzmsSt5fULYXF2mk37GNtbcFuB
4he20kME2ACtizPhEzsr+dQtb2ySo04VLh3FVB4ZBq1/aE2JI1Rx2Nk7zqXkR3AnF9HvO1LbwuvY
3QyQkXvZiIxlg3gAwXwTcCmhEL5qUdzkne+FGwq+uYzIrHVaUUFA1UVgDKa8ES/YhoheEMIRfzxK
hu1XM//TcxkftqD3YD4mW81QWe87sD0EgAxbMeJRfQv5DKdPSQPoIObUT7KZUkyiNh0mEimCQkqx
yD+YvGHvJZyuYR5W77tTPiKcqB2xmf9981tFwUwQh08kBR7ySRac5FPXMD7uAzH8fcTH95Iffafr
pJt0na/5BbtlK+nTPGjFX5h6Q/yH9keQTLf44qgg6NevJ8JcwMSPvgS6a8IRHSYQgCspxStU2HoU
IBnoM9fux7E1g4VOvaQCXqslKHN1eH1t71JqhKzRUKIjvNhkLDDg0WqOfYpYNFoyxSRZxDT4+wCx
11fkvS2EC2TGrozIndf6aourRWfzDYOBjD6qPNhTBWDFPPoaZ33z+iGtSv/7KDMQ2+DhQaAYc7wB
+VgxO0+L9vNMtcnFm7kO53zW1BUaarc0LNAFVw5hgjs+QdItfZLoXCU57l24TXe31bPuuDIvG6x9
iCyFgB+FDNiZd2YQGLt+uoTqi8GzfWyJFDWcfBSCCgZg1OHE7uxHGlRfjAB2f2wjcBnPMIlDlEZ9
vaT+yhdRSGilgriFANkA8JWD6jZKRxuOk1YgCV3HuWc+tQVRSL3ElUSMHu7UzgHBClK8y1xfyU6N
AVSbU19NxyLOKaoslHOa0oGk+DYyom57pKJHBLwNKbcc56QQ14eP5yD9t5xkDb9bAPlfzVP8bnT4
fCu+dCHrZ+blxu0nHiftdUz6TVybHVy2LctiiITMjae10fHydKHRaN2GRqAt3KvMl8NyUq1H9EAb
ATRlfWgY7hcSBCagDIkCGYNGqUxdMCY3dOvj9WJvakGtyXCh7KRQZG+OXUN+dJpbHu6OrUbRQBez
K09kVazfT51qUIFFZozP25ZhV721nNWohQy5DeQ2FEq0wBSW+8w8ffG5UNhl/4BS1e7I1DBzkNYP
PzsNBoxkuzH9C7hAwcvCI+fVuiNUbnI56Ts8Y8zX4n2kgiP8JoN5GudJn8SPHq8T0wZZhIlVLTp/
y+/4sysXj6xABUJ72rfS7BBrnZxftEpmM2U8s5QNdBHf6Fpw86KvGZ6ELKY0C5d4dmpNxAIEL+hD
qwZq2qn6AIYMb7VNyOkHgMfLrcliWQtp2peRxzFNaP9LEA8MPuX6193hWnWeb0d45RL/fgL4Dpeb
eLMU+jBXcYyMxBpfPWTHeINnrtnKcCtYBi50IYIe1YGym9qEt5v2o0PyJUAw/661ZE4DJDIuVg+L
ZrYJZw4nIko0CaT0weOlUz83PLh2u7cvbEHTBJsPi08KFDNE9fSzi7NRiqwiRP+KTW9uVfZsSaPu
jDZzg9x2is9vnQJmt6NOYxd/qwcg65mmm3s2NWSCITk3XtWpFubetT1vXew4GdvXoLabyLs6XTPj
mESzWViyAfBp00bHDPF4sryM3ebb5JWb/M7TwbGtt5JBixJcCeSSgulB3ad5V2xDrqBe6IigC5Vw
ZBDcae4Ra46mTaNHIhUHqRFrxyRBEMcnroOpOBITIbUShvOQeIyoFdD1gYRS1ZA0RcMt10EF2sWd
zdjC41qk/e3wfao6ywGCygfvkQc9Lzp3YAqRUQ6nIpdteVDHA7YkOU5VPCKzzQqSbY1U4yZJ0DeO
Te8ZXATJRJG+uRQeZ1cTbPCaQ/bwsedpC1HHplfGgfeOuILfAE+V9dzoMXu9jxR5hIcpCfLvF1GO
5CrJDDnU0iT0RsBmAbzIcLUhxICfhpoNgoYvA/URl6AG8rmfyhJFZm3mxfIEThGDm2/Y/CnQ+hdO
GNgO89K0EzZPDfO9KhsFta11LWAzjozqlGOcPXs0LYAOU24zZYGYxD6ZnBn8ulXsabuS4KbznFRd
rhz62sRVNbfhDTbe7880WHvfF2nh2gHcPh2b19pT3OUuhl0i0QttdZkUibzq0ZJGYs3wehoUbWqF
xkZcpS3cmGSGDwVIQbLUBN6z+eFLsGfAFF0ffZj7xaNNlha1q1LU0hZgPf4qMfMsjJW5squksod5
m6hgZ4LN0h8C2+rk7NJe0uqcu0g3t6xqlhg7gAuQe3VdobhnoRElYTn0Hx4VP3w3ioZYdca/BGJW
78AGDoExPdU7P+uiR/zIUmk9/TXaFsuj8+Tx6wdW232de2A77P0ikbQSw3nBgDHSgJDmbRjc+Y7u
5n6PjO6oBnjbF4q9BXrnGdc1Gh6WUUvfGBuiTkyiGQEbYdocyo2EdU3N3zBRi7XtImEuQv05ZtqD
KBDxMgniXDZq86ibyR37bYNDpJMl/eS2RQfxzIcdcQxzFhBt/quQcRWho3rQJtg2gqhdHGFJZMCh
YWHMcDbd9JnjI8IHMcik2XjvSxwmnvtj6DtJ6YyGlfC/refeM1HIr6pJeJBUZG0zat2UUC1Tnlr1
ib/aWT8Xc39UirFAh/KOUi02Jm1kHWR9RUITKK26vcV3YzTf41wbE74qZ3jE5i77ufQU8c4bFliY
Jx0WVgN9+/yfCvpCnH4HFoS+uVa3vMJH8JZwjrg1TKRx3V9UNcm59Gnzkpvk0BkPS/hvABusAXe+
19tEOoVaIQaeELS+Kl5KMCrHoK931rK67LD+HyI1hf3gnj2wpUeh4hFYAeHDCZ/MRH2a7vHrt4Nz
xK2V1RtRHfcTSgZ+1MK+wWbrPR3q0eqKCkEPuyVRoJG4lF/+HEJxsxWp9sFjjFbQEHPIkC0M6RLB
sKpoNNqQ0gJX0cF254MHoN4LstuFoVqPaP8slPWFHHx3uDNlJC2VO6xss0AbCCL0YuxqzIiOld+J
s9JZoI+b6wl66P3etiq4BMLgBhPvXcEqL9LiDn83KDGATlAT2ydTckwXu77JjtTz2o3HxqK2q12a
gjG00MZmf+ZcrsThZDWAUb5yBMpDGQnXun76ccbEOPA774o1h4RmMPAJ5C6gesGWNh6OqLze8Lon
EV9Q+X3bvpPRGpOTKI4/gdm5GvVY471CtaEQQUdGpvZ1fqOJgniZo2w3VipUXPGAmC1NqQyl9Hjh
41h7J84nz0pVJ6Kc2/3XeIJTYIDV+fe8TiAcdcoHiNo42onp24WYruclyrFzeo7bs1AS0nfKnyFg
GbwGBkwbztNCo4oqTWd0bKO/L48rCu52lmbLskA8UWCMvvAe1l1FVVSF0NQ14nkLH2hCHVwhRUSr
Jw+Of+RZYzVPoGOE2qA6PPHvMV+ERTW68bzZdtOkU/bQeWqqw5lOCcZ5qMmfm0yLiDmgN1pWnfok
5XO70g4brEJqDyEeyZR5BbCnWTCnJqBpthNJatyZDprFeMBV3UaajQPzU1PWPE078Ntf11AsqtZB
NdFfHL/db8ksqOsm004PNTVI98uRYegtZv4x9SxM7k9C+gWrru1zvMEamTO+lFzuz+9ErJKyW5z0
eYgLt0G/If4JhpPbZOGGeZ1lzDS/shPvzSoxMh/xEOePWQWlo6Pd5fu1wv9QU/jSRHNTZO1BoMi+
K8QvU3wzcEi/nB61QDJLqHLWPVek98Dq6EjUhKMgj22ZeW21zJ1qYlw+MhmYGFm0Hhv1sNTNDCFN
mkQVic1dPufspfEFpbwjhS7Yia2AJZKMeP5/+2UtHw0zqg4xpI9UCcOyqd5Tum/i1JS0dKhH0mrk
zydMLB9tDbU4TA1aCyrTv0VxXYsLBOCkKObYWflcfNef5LtySoD9GlLaVeetSjUa5dt9Qe9JtovG
koC+B1T2ZuRMop2HBQ+y154zeusdMpG09lD/FVb9gdW7qB+56G/FWcRjkPY8qMb3xfDfeCdD7cA6
xDt1gHaU5EzD1N9J/lzZIJF9L3A0wQ/sS9/pR9aRcKtS6ABJQKp5VyE54M4f4bp8iG+IWMTAwPPE
ZoLZxa54ShGpWTNd4KKI1bQrL4bxRYkpDKTyU2cfdjdy5rwn3cGTiKhAkPNgeHbeg8wvIc6Mwu6Y
jITc8ry675OM8I51nfMMaaLmx5ukLoMeW+tOHO+UAlrbB0w2oCQEGa6UZvR33ssyDK44l9j/hlWg
xmpgzVLb9Pw4U6UeLEaL7vtTxcNEGhe7IqONZhaXmYnwwDMmlODdTJvEEcrpROU9YKwn8v2TXX5D
5V4gFJ3hYFcvVwn5Ty32lnbRUKH71vXJtdIVYqN8AipuzooA0fchcg5sBGyNBTH8bh188jqLW6lY
qMMq7KoVITC1mKJbP1mkHJUA9DEejV1oCY6vd6jK7FaspEpO+HpNNQ+OlTZgYfnlVWwsXv68oe+4
nMINM4eE1ctBZrZJq/BQfNfUJX1e4+KbnE2ii7A2cBL1Yoy4onzCjMhy/LqDRFpbgqwmxN/r+Yhr
toARFvZAscbw6IEeQk3lU4gVMOti5LiqkooosWJtpgu7nUG7PtHSrT/ihI+D33lO1BpwD3sclRoC
RMOLvYuw6oB4fXikVoPlv167VaF+XtIpsztHfchGbT1g2+biGuKLsMOQ/swYzFXV46XCOBf+etAi
ZtlBG9NCLo1BsNcVxdtVXLbFjlDE98SHJ3s96aPvcGMbMkZT6nxndAZeMUdntBK6d+pALmCyROOQ
eKHjOsMX40A5Nez2MIYll7OY0lruB2OabrlVakR5st1mjQfPlheQZUG/ThfQX4RQkx/xv0RyJWHD
85izY8FuVJkijE9oE8rJtJDFWcIxderZGSSoYZnq7FlRjCIHt96BR6vDR7iEQzNpLj1A6srrzbke
mnRq4agJ1V/OFDPgIJExvM01dtwV/sW2iDUz+DUp78ReX0jx+ywvWOUMC7250aZf1kgv3NBd0bj9
HIkDwVJBtYgNKruy0dNx7jdPt7g2c/e5BTqAPdrdXi1OhsMcDdwMxz/YdwkSROBTcR7YyxYk6oKC
6shRkps0LMPPwMfFWn1zuqJU8oqe+AdNe0F8XIt5sdYzAJnKMQrPilomyL42/WfW9vZAvHSxipIr
IS9qhPK2/gt5WdGiNqLBUmldcPyfl5bg/JdJilFmnuM9HSMZOyh0yczUKvB7fUeQ4B2IKe4/JucA
OVINL629ZRytmjNxMHrUXFbPwJbID2k0Ty9uKBI4C5/I9aqfqZAbyu/UYLisPX/RZqLbNgwpD3Q0
wJUVd60keHAqIvPOyLRJF+RshyAc6U5dkUoqGs8C8Qe257yVGScvowddnoqysC54DXt6XyxM8LiH
sqK5dOR+oGMYRl6VGSXDMTdh6Aa3MwTQKnfL7E82IkxocHnAclPT3Z4uUH6MTCKRHwE5vIbSFqOj
XlSoSaxthG9BRg1uzT2NckuHmte8fn/pAw1PGp97+/NCQhrpWqEv4LWURZ4NHzFy4XTgdKqCtSqZ
pN/1V490ZHhL8GIxkcAc57XrINvcTxM9KPTqdtbTTHZUMN36xntuioEU5IVgqljYZ4g9/W+va9b3
0DDSqScyR3LsQJnVXIKejGTYOCVmksV+CD1uJT/R1msn8bUKW8ubHuI/vRqDTdgAO7/tCW81ZiNA
cLEa16K/vCRmHab5bD1ev4n1o+Uc4OQKDfvbRZ2FrD2AP24e2piYTimuE2G9dSgntCnxDMFVO5ID
LJKDNjxZFav1GGY+3c18AtV3ne4XH7Kj9xmztugNpYE6TsaKqj6/8Lqx5XQYrKBrStoxITjMeskv
e2jUgCeUj+fJA3Oupw8Jgc1WAq8I0poL3zr0TfsAFjVxIOPrxpNU01wXV/b/ab+L9pEtNiYlMqFD
Ev2L3w6RCSquvCFG9O2fb4Hyx6dfcuuipk+i5Yo/UW4YBf5qETuccm0DCvrJkVx9zQRfKKZeb9S0
A1a9yanrlAywamXtBnJsiDpkOsPa1ozcx+hWfHwYG6eKiCHsGoaT/mID8sG0ScSfPtbuYtOa20Zd
+sPHF8PUpeoKAe5y63EETO+/bR2lTy5BXOfkx51dvL4WkjsqCYGZy+4nTVhYGzvwkiqvSWdCHjm/
bAyLR/O5ByS1ipujLDNWqNSOnFUeCOydYX+KqEUM+wLfOxQy2AjVnOXGx3++KWTzv3XLNyFBUpia
lV/Sp7f29IuaCeiOS6UGXDfxHtweRXeHxtA4dl8e+pz3+P99SOnninta8vvGqxYOTc6T1+uza0cR
FYjMHcYU6Ux683PvTF6plCfss2vNhTOdMuC5CtaQROFbMscTIib38rV48nQ9mUCI9w+L0oCLLWRD
83mr4fn4F4OL2Z7hhH7TBhxLcrnRP1EpLZjJ8KfylnJGUl73m431LTtg8+xDdW5/6p4ANl+7rVxM
MkX5sFRfMbVq0ZfiIRl12oyi9ybT7zTLCILNjxZoF/3mU5e0ZWI00WZ3MJkFHyi1dGnbi2x9xfmR
xqqLczpt7xHa3bMFMn2F63uXuu2vK4KOgKkRt1FWhGyRrMZUvnnSsWoKN2XoEWwtItrvDpbeI9eD
frAJDWe+xa6AvGfnxYxYbURou0lzaSoOwtst6CJoMMTFrzmyiW64NRGz1illFmO0DQ5XuFVuAp4m
0MZRtYL2T2rvpnqkws15065SNajn1B7Ro9LDRzOEGVfyp7+W0EMtBAGl1aFDtOLqihdEzEtPb685
GRk+KrJHSGm0EIJk8eGWz6tDSkkD+6bYUV3SCDX8pqOnBWQtC4ANpY6pPlY/J0/hWTg1qNEKWlQy
cOFBHAM4mNjro/ikXA55g5zZod5TMGlJdawJdtjX+SRomrM9azUhMuSF1Joz1jQOtz7gq1XofzxX
stIvjnL7Dv1d7CKbNY4tmDcGrXFKQmJ00tB+tlP7JLxTCx4PH8zU7Wy2jNuk3yFlTXhl9YSpPekr
X9uvN9usm/n7h//ole/mUSeKiaebLsPjE5VZt4rIWhpWDXMizPXReEAo73cmFlWtRO5qOlqiu9is
iJVwAkOQ32sF/laO1iIzyccPjuwANKVTU2XOPmfkJE5sdoiLA8cT9EGgFCA/2r0rW7LtQrLM8oRz
ezB2/sf0s2zCNoZ6dp3/llN7u+pR2TLksHYh7+LdTKDkPNUDrjXCBArQHeIY6tccmkHzoY0jBSnA
av4/L8t6iZ+jHO1qz7Uuq+Q2V17eX6j6CWJFycsL0+V37O57tcw8GEHOtX3D/9SaZkU+D5dz2n7G
SvHzKOlshz2PEiMsH4Fs7ZDUAhbf2mGECvdS0RsXFVrtbDY3DFISWYGXItV+TpgIIk6MgLUO+LWU
g3XcTLSz+azPE0eTbMTGYYyLBNKMzzhdxKlct7V4krVS+4OUvHIolq8t29BnlCNqmi8hJXVlhJs8
4gpyqEQJgd+8DgvgK9lWh/aJr9e6mlctvy9wYYMo0fhMgSsBLH16fMxFYhAfEV37Nt4GRnTL1enA
RwnpqZafMJBy2eZ6asALSlhKzxNqJ4zF3BEC1VSiEMNVFNV1HVroEkHPSXnKEZiG3DH3YwSUN/TU
/v6fb+g0X52KJkpclfYrE43BywZmyvtV9VdfrS6oLRdMuYtwm6ppLUc1qcYZi9U2315yTB14ZYRT
R0RZOvyT+GTeXiGafnF9cXjUFLs/SnGsVB0jteskcvoZV9CPnfGgvOyfemPYNiNL1LG+CsE+wpkS
YEKViFYI+8SGbrFthVE+PswWpAuc3jF/W0ALTA69rBkHqir2BJuj09RolSqK6/9AvF1sVN8cYde+
7GDd/vBanF+GWOVhGItJh6Y2z/hKyd91QHEl+TUcNNWCLeggb6d7vjngpgiPUHjFkRDSa/nR8Z/d
yo5vdFwT2bQYuTARGWsRODTKkWKKldrjudKDIfC22EUhZ4TYKHukTT7TwKqbp6EhMC+nyelhWQCA
czajcw6Z432Gr35alXKiwd1R52GsCTYWMFkUbi+0T3bObW31f2xp4dwTzz9uQHD0SXfmfh4/YfsF
Qa0p0N9GFvCybtKGKX/DodULuJ10dAJccSNsEzQzfkidtM7+hwYAChG35hrwoNSU4DX05ecaBTOZ
gbJprK0tCLDqBPPTI825LrwhAftrEyshPFwvn3UBHx5QpZRvk9xNeCBJVcorz3MMeVU9Qd4JAHhd
bshipdTdGUyassRJFxwMwDZoVEDuF0f+5JETQMh+cP+l++tdWk6FF5+s4BXK9qL1b7bBHzyctGBv
/lfHsCTMuGU80nIiH70LMQh/+tqk4VqMBvarqWxrdSW5GBaarwI5QGnpWU78DzUem5IJuvhxIIQ8
1FBL21JpkLBbW0XUUJgF2YnvaeLktW62uEQj6cTW7wZO8h8LJBW8UuoREi2z4tq7RXothOXPAyPh
K/CsiWa8y0Q/Q0o2lXmUbQRQozTYESRK4kft35qMruicpEhbGR6LEvoyUotFfJVLY2YH1kYCVMa1
ehHd/eknLGScsK2hN/SNAaHIEmD7ha000DfUZM8ZkEFBDu0RhKVO8VJTVu4Strrwlp+GuTgMCLGa
JdS20IDis8r/uzs1RtBJObCzEKJCFki5GAJvZDhhmHMNY6nRiqCoIuUq7iulXD94Volc1fn4y7dB
dNqZv/dxPLF4dAtRnT/Sy1MYB0sAS147QHbrHMqfPcOeCFQOekUPYYJEffITIYh6G2HdrzR6wKis
l8bGbAyAs67pLNMKdxX1EM1JmX3jRchjELCKKgBeo7+kQHxyK5B1Zn/EibA0oeN2cDpe+MSIwSfc
OJ0Zto+d4b85IJN2UB7Uxce1R2dko0x1MkisfTeFheO8PgUn9ICLZCAlM7mYZ4YgzCL6wxREbQ8f
pRXLbqIO7vJvk1yTaUUnAVjQbbY1EOJ5ZxZUh/k8g5MaVVbTyRLAawlOEN21a8hTsfzbGPXAMRUn
fe9Ptvurs3U9cySn+Z0NGz2a8JU44CIR+1sXe2/xnVX7dv+7efGbxuM3J2Hj5+Bvkwp++nIACKnc
6XHiQ9wtY/txjlLZ2d2LhzjceiskuBtaBdOBWPuVJ/+FzT4tAjTTG8H1FRHRahnZpMG1cCYEpUlG
rqcHhr9jLEtDjWEjGmUcS9sb6fOfGvmyrLSM8iTlai52zGHH///EpKQvYbymG0Hh2fwzyqSMNaX8
g5yx7+GGavfdoMVhjm3nuP6N29potS3mC6MxxxiXpgmOxHSohb9EeAo88zQhdopNmWqheeR5EJ5V
r1h0DKFnF+z6H0U6iV9S2UEnZaGoZkOqdqhM/mxCE/YW/0QSXILfigwmFpa1su0J8XfoS9wkHyR6
O52/m2bKPGh76qpkOmFslXnzqiqCcl6rn6FioTzIk+bqwaVmtzqI62PK8pU6ufauwmZM3f/zJxPL
NrJwegaQBAqDq3UoBsLPdrPtsdWBlH/ZSoX/bUCiLZ9W8o8G+KUPHDHIcyxcpA2u+qxcCbkE+aBU
wF5M9297TCNK28NBx0tcAtA5skd1RmDOtFRGJLaY3tfj1kKJPnmDQ6UkrsJgq4vEyU/cIX3p+GKn
7GZkwxRH3Xpgurv8oHxnIQ/hcOVGK1R4YhXTOtIbp4HI+KxyDUNRPJerOEtRpFziPrHxavCVX653
EYj2N4em8tqVnb83YP5bQKpAp7o6PQC++MqrWUblhfrTS52+HruJtkOTWwJQDFMIMDUgy42t9Dm0
fwBVmvrnZvkURMVLzSS/9P6YFluhZKC0GiqDrmJeVP6U1WXrosIgnBLGXtd3xvWo/ySOoAGgXwbM
EfSPZZQRyfhwrxky/bp8yykKw732RuTqwJhOHpSFeqrLl5DDJ9BC8wYvluUy9OUzeO0u2+aJv6LZ
RcqaJ7MjBYBmhpzHiRJmlQdbxwT67VaAUVk/LqbLxUvwjYNZ14UhYwOhj6QEAoUXrD0QislJq5zy
OrLr0of6NA7U/as9VlIq00OmC20IfZ30U7ENQvYPQSWb4cL4enzoNHFDljOkVgjfMT2YQvrtup7B
rRVofoi+uGUL9NGmr5F7/um9igOgMCMp2Vlh78qNWaumdNJNEvyLWQQABZRo+p/a2bXzqz0XNwiN
Ec7ZCnIYmxKKOaEIvPAxMCMSwH8fHYIJpHvxEJNBAtU4kW7MldETB394LDP4KXgBCo8yzwHfRXvs
zvoSxGZj46GfBkvlF+Q3eHexPPPKtWqZfup7mug6b/fHDTdPVgYtId3W3LiMTx4V6optgWR4axWC
4ogHUWio2RHStdpCwNB3t5xOg1aoSVT/XbpocG1Bj9JqwIns2ak23/Dx1nalytAaFRzrFL/6GvNJ
vTULaons96AX73MzUjeLJcdVJyKn7raRDqamMHF/xnz8O98AlVL1y5NyV8AOHTV2B90tBxJqBQTV
sbTzLS/xCZGMJ930Vi/D7zRnn20ijlsrDuk7LiGscw/esaYeluhbogdx57MefmpIM22IjsiiUPWC
oX1S5K/hrnAqaZXKNs9IDvssNwoK1mBFZ6si4cGlmPSlqR3B0l4agG/g96Xtvo/37i0/2W++BYNm
HhN3gfVv0GKoPjf9vcm2lM7Ljknnj0bk60xDV368tXPx38wUhvHOCN06467TwT8Zp6nVfvCocyOC
t5qPZgd2zNewpsmS4/ILeNSi4WVtHnjB1vAQdgoOUCW72M8BzedbHSZUX6DpyN+q5njITSo+kNXE
+IlNrygsa2naDlzHI/ANOUZyxRJrFlN5nLAIw1u7YwDfPyr+6wmd6BzbsWX561NjND8QH+nojxKt
iaB8aDEJYMVuv8blUwdHHKhxbuZSNUep3bZ1dXmGc0mjUCiGS5Ld3SSRuqh4tRY3EUrOtAzwH0o5
76qWVL9Rpk08DgPbFWRfqEn/1YjuTujVKCW5XFCTok8l2z3oSY7MpFRDWcJIrRL8np/wC2Ev8NWy
+JzxWTQfynJ9JW9Kzq2ERysKTAnssQAPpJC1VUYTyETn3NONJHIcaeEe3vyXaJKAuZSjALageRK4
VQhQKZx8AdCEy4fDaHOeQZ9DlAKy5aSW9PK0rT5DlDPlNuCB9f9M8nGckVq3qbbYzNnweHUHpf5r
DUC2hj16ntzKwul7Wgo3c3ZsfaBBRnrHpQbMGFKdKUmWOkqhoY2x+msYkQUAgEBiD5LiulDzSRZC
qDaZC43T7y9z1wyTHPM5ppIRg/R1ceiWQRTJx2mKR135PMXHTcLPp2yN7jMbZL+CC0Ntn1zmyapA
TCe6D2MSK4J5+1gfC4tRvwpMlwj8xGGlyR9A6KmaYStb3az2f8gifwMYDVaQRPpL5/lpUIYRe4IV
2VCRnN7wvBEV30NCDL6w76OX/rfqY545otfuy30vENseEJnLYnaDZthsWOHvOa00cDRs2MatBARN
/YvBY0TbiuzLc410nJ7QCvxlohV7QMhaY9+dUPMln7EKpBbGqgIvujNtk9skw/Z9taWzjfVKEVhw
ynSOfMeJ9KlNQ3KPCvKu45GP8PeUNOpN3B0PqqYW6BNjTQcCjAbVt65sSytDDvh7hsH23E5LMQKn
aipBidyIl/K2boVvbWhLb6A4wugKtZFjGOfE2pW4cqe+F+j/x659tWzjk1XWLvgHUnl2pPCfYJ2I
Wqax43YScSSo75duyZJXKwkxKBncV3g+i2fkOQrsz8IbeeQocVm0hA7gdv/prMYQas29+HPGuZ2X
Dg4vfWOCXvNvZyX4Q3MTU65FNdneB7K+EES9OnnCdWKnQk5+npXloYOageLN3U7ohe0S20VvGoEj
kELevHHfUghVXgSbUSHhD6l9I0kBiSs1Bs0H2uV8OTUjMgjZvKtakdBOw0sEwxFsKOb/Y4PNxeML
KR548WLTBuYeJThRXg147ReUTdPADTbXPZPXFsT8FakmpJcGUCERneCBzkIe3hvtPSUl1YKiaYsk
IiU2v68/cl3MFyJYjVIQU6CuI20PghSV5O54+Gn3mcEp8jo9e8adWRUrUcy+VsC+SkbJ3dNt6acx
3AroiLqmxxTRG4e/NwEyTWdJyKBR+RxUHkJXCz+uk2/xI2iZztOnza21kaWUVHc0+cOwV43hI1pm
Wp3kdM8T+X7Unfgr1PQ2zy7wn1bEmHj+5gsDe9ylqr21WZggHU4pZ0mI6zXcMcl3BN00tWWyvugQ
8cW2irbAvVwgpzKmZ0TtP5Cbn+T8OaLNIqMxlYSuXBn+kIA36rTcg1XQHMjAQ0y65A7V8+DTOA0B
IvDeh3O/1lxDZitjr0v0VG5fwKaMFmPXxnz41w85wYfVQD/78D0qs5jj0tjEKhI/3IS0QuUohwXU
xnReaXatMt1j67F3yn2F0MDk5mZMM1RNPXHtB4BmZFaTYorhXUG0I+Yho80JyVGP5l0BAtBPzSps
BcDVM83wIqAN0n94v/XLJR1SZz9mQkQW8jFyKpKP+D36XqUoqLPfHGowWG1dZI3fD8riYphj/g8R
RIRZkgBSi/fSe44qr+zYtMPkRi6XoAlnsbtcGTuRTNlP+GqZISK31ByX64e6Dh2W9BT/xMUd2k06
BvzEUOmgQxo2g0NE2vud3C3AvExZZvXbj+6qKQc5CH8H81kut1NzryIQGu5W7QxZcYCgqoMDP66E
kEXjeAtDfdiSs0H/frd6iY5ULQjWkxZUrpZXCNcbpxMiUGMsIaI5HyWzMh1DphzdoZNDArQ7+Ol7
/mQIc+xyLFGA7K1Pt0lEjz6ke+evlqnVmDAERKRlcxqTPwcEXi2XGlJGsZGBVylHYTPc0Hpe38fY
WQoVFczWOL0oK6eGEtBVx7+KKDOBzVb9t33+8q0uvzZ2ytkn7/fDCSEd9nqaAdDTO2DGFTJolbwf
l2WGtdGfJnbSg6QRAzqfQheGoyf4gGppbX7YYaAnE19wFK1AC89c6YfzSTIQ2xsCv4QwSaQOUOzC
zqTc1ScBuuAhm9HgzJNAbE1LDMmwza1iXK+mvz9w5vJoCajyEJ26lrxUjd/EtzbpvhqHV9cZvWT/
dT/6k7f/n3iM9NhwomceHtPNwlK7C0J09jzRtQPRsWEENASuc0UFpaneOb2OYuNy5UasYh5KuWl/
D7NTBHxwt2+Byu3nii3iiHSsi1oUxPIco82qnu625o39dHnqPoF72NSqScS0pYaYL+YXMiDjs90s
x50g4YrCoDknxugh71wEw3UqZCXl9aJ46+AjrzKVqSL1HSUPYcH5Elx4DcUCUDs6pHOUloWCsPgk
pJfLvuJ1UDYgQvoZqfIsD6p+010XDfViowD6A8E7XA1HtUNeyff109c+3cKy+/W7kHGQZPxFHYaG
/IYlbTw1EWkHQAbR8oMp+3VamdoYh4pmtaw5SVkbj7894olJ+VL7bT95yrHgXNNEMmBrcwUCEFqb
vOhbyKhY3I1fBffpL+8BgLit/KF7ft7Bq753Fg7o3jX+3ZezUwpXQrbTPAgNubiBSlIPYEejQEfc
u9+mG0qfBcUJue319KA342JxvxpVIRyphGvXqdiElswZ0TuJBXLaEtzf7frJ+qz/zMDHEK/COhBa
xRItyO3b1odlmT/j+ZpKRAqPGWE+llEXez3WV86QAMUoBgcss/I9ioB+0O2tdOf80u6C9MwS4uBl
YkrFqbaw238L8JoRUJ7z/4V1qgivVuZSKySLCCoc1j8u1/tKTisKUipFD8QEiqifoH/ZU1gQMMvs
41S22m911+RbRco+4soTkeag0zKecWxEvhbk5XPjJ5MlI8gnpBahQJDq/uWLlMjUGwRF+CYv5xrH
qpS1ZoHK/qh3EADtlFNDCOD5Snfmnftr5dMBGLVRBZwqZy0fap9XNAFSyNciGLmNrjqfI2xvYVgB
GVZNbzghk6agUdMj2vlT7EfBN4CDvY4VrptDdDzsNuEmQP4YzYd4nRkWFiQuEVxUeZMrU3Ck5MSB
P16yCgbY89s9shGwcszLiinTKGUPkLjYdSdv7NcK7OqTy2FMkI54GGn7bT+AbxGIcZcYe6ps3dsc
eQF2ccQtorLPOYDngXTwMHhsSh2uj+MTUOSOpg8Se99ng0rp/plHGpA9sqK28F5sQ21qfDtb/RHN
/PMJ1Zcx7m9fIDWnbHTicdst3+hJL6qs443dnw55lxhupcAA33JMSKfq/gqNVesw0ZbpdOaidhUU
FRf3MphHjX8esIOt7JRUrKsx76prYP/ltv+u3uu89X3GD2PzESJFFySCu9RJlW2tbEAaYQfwWXp3
uXpmB+vPJG51R5jSPcFlWPw935D+6AFURsiwMkUuLFSooBmsgXn5exqP97EB3BEKmthtqZ3paNwp
7vFxqxjibF+7I6qrFgRbnizPh0RkQnr5jR9zgmiNEt4uY6Wdsw7LTNlZXrueklLgC3PKqZUP3nca
r2RD3IANc+ow61R9QnvcTGQamab5+UY6pwxO+Y0VAwyiNoTVLTyDWlGVpTftKQh75rlhWg8CO6xF
DsSRD0pa7jOE0kCrNGX20iBbfRKh7bzzgTsMjpF49lh7sRyqioKqOp4QU/vac7vLRR0LIJgFZ7N0
Kn80a+Fz7jBGC8L9NN2r1taClScU9Gnq4rU2YFjmptWOlRwaipc7jtoG1wlAUo/qoXh3P2zU4pAE
TJd7683EVXdE1IWGAfVer4fM1Lhl0zsFTqcEq7xGNCeWZWniS/9BjnYELDAFMeEwBXh8Q9ka2F9k
1SEYG4jxuoiKd3hakr07787HCuJNqolY45biWY7UgvLlGbuYB64kIO+yUk6viAZxDPpGzJpDks+M
I3E++GTreh+QYTLEATe0ExCD89UJn7WOf4wPT6n1qpSicMyhr3i9k5h2H1kCAQiz9YH2yqfept9Y
n+EyuAlsJ+VxZTjYaQWUXzc36EEoxhiLJD90kK2P4J15J/oxSA36F2+UII7ZjaR4kcmixeyZbT63
NJ9PXzVC3VJLQaJ99pCnqs8mMSBlad3PePKT8S3hmiWvXCtybNTCamKRrSUBuAwr98QN0JPpI2I+
OE0GEPPTDO2V5Ok1QaYq4PZAtTd7R+FLHb40RzIinzEBnysuuZbMQp1kqMaIi/eTWA6YHDaDKq18
MWQyXcZYByGWFLp1sB+bfw/CerFIfL4y+6b7fy58kFZaWm9OI7J/IhXynPNg7mCQVr4Gl/U+57xm
DCtXgqq8eAEKTAYIF8aYaQp9JAyUSAYRktHOMyivCX4r4UhyuJZ3dDyjAFMOCJcDv62nSnizKtOo
hD3y8y3bk9BpgEQPUAF5SSVHTdlkV8G4ua2fpRU6BItjBnobBCV8pP4RpAWcH1zXIym232QQhW5y
cnvrQkNM7H3psN6hyqnWiQb/HSzXj1V7dWB9ADYDUm9Tv1aXrSp/BcWviFGFLdp+7XpSBhBDb6RW
m0ElJ8t2WmFIQkZRoUAbsJqepSPBaQvtPlU2FPPNwmBffD/3cYgs6UvyNsojui0Cc9xaIMlu7/G5
QfxSECyGfe1u7W3LgcXs94JwpZLBb3GSqV/CNnsAKOLpyYZsNLKTzV3Lq12qu+e5RlWP4JAjm5wc
fQb1pA/4RSO4iwTI/NLwwA5ZI6LxAOfC3m9zAQv3vKPdiV/iZ2CKTkUUlgr3Al0lg8GQByfwbf2G
xKlbv+/F/+hKdWLSxnYshB1xy9sfLHv81aifJ+w7DpNd528B2P0AnxCYyRyHJ/aC+GBwa5IkQV5H
ZsJS4R+xgONSQOLQNuvXfQEbXrLCUBTua85sxA5KLbSXFYBpOBRJXPJ20lNmkBc/6j1w/Ixb+GRK
qS3uRtrPWzg01sDsfPn2ghj/+Mk+YlEFz7QQRt5KNiyxUAzJpRdQdVJuMMio0aMbRxXogyqXxmYT
VdUL7Ka6FbXzSpIE6fZzW+bt2I0SdIQ5R+TkzblW/p3iIH1p0G5vFPsssjvVPb4R6pON4raN72Rp
Oin2NX93Suh96r+vSiVmyV7+oj1shwUCkw9lkR9YGtVa/im9goRwN002h4dDl6OlqwHe/5+7YWV5
LMKKSfiRJnMj1ZjMjMBsZASRIkNikEsNWgCjYvvYYEls5k7TTmRBwbxs+ESmlFMu3SsYCUl+3J9Z
RmFwnAqTgGhRcqfF6gf9fIluVmYGWLSjwQOVFFQth57Zil20aDVchfQ0RavVW4aVI4SuS4gfcJ2O
iqkR6qc5LMVSKqFfVn8C0qYzRY66woBgF8+kLDTojZ7u2JSl9DibwKHZ/2vaueRpJk38fa72EJRj
zwDkT8tJcyehBzkF5NHtZbfagdcxPJ7tNAd4Wsb2swm9X3sbhphMN87IlhVmiHuFAtwgNtC2i1C0
svNXOELTDvKCdnLRcE14Bnm2FuHony+g8wVqM00RahKmkQmZeIbguR4E20rG9eUml9n3Ri6lXB89
oJjBKzGxCeTrG7nZzimz/XksSOXTKOyy4ENcdN+NzXqdf0NVA7aSUUBF+nnqOGtsrkrsBnqkrlFi
5xkifTFXaWnVc2H8LNK/Cuu7KdT95b1DRK6kuezatwYvuhXFKEc50T6E1kJWmmXjDQOnkVfURnid
rlmVA+OZuCq/CoJOG+1fEtZ3omKeorLfsMUeCMEZ4cd2KCjorZoW0JtIn8n4P2tMhS8sUhgNRr4n
79MXLda65i60Rd/TsvPJ3qKYLlasixvfjP6NtqjAn8fV6EGlVZF8uj7SU8GOE+iXuCiB/tjB1c2z
GGbuAgtGDLK4oILsoqbeC9ozsKLx7Zt3abTK9f/sJvVL3u8aa2YHT5pjKizLjZSF8SmNvC6eVMws
7EA2vsvsXzm0r1mDZ+c1RjMoet29zd4Yf/QZWBXmOXl0hVcZQl6i81GjcHkeShI74z0pn91GNiNH
Y0zEggZ+u5OPNn/c2G0PfGVhFmD3IaiwlZkYsVEP/9gd4IBtpffQrrwIUyHoRU/DbO4LJrGWkn1q
aJIx0MZu7aOrflV6vcu8GsmIfC6PiGmUuVL+ww8GgY5LyKnlOd+Qjmf+K/NZmsz6SMc+XOYZqjwu
oGXNJFtJji9rb4pCMTOS7aJh1jGRdbmZPo37HUC2KsT6XJCHo3CI48f64RSvql279ab5KmnOfBIs
FkeiNtHVquRpMqNlPYEvBXVynwvJGWV6x7ZbrWatIOKguK4wg2odvXK60v2Uhd6W6yW6GLTZMU/9
ysIhMOYZ/ULfd9XMjWSysxOFkbtYD4p2kinUB5XtNp3iG4edVoMLTDeiYWC2Qw89d8tt0qx6YCqv
SQ5fGtYwYEHrKWaTB89h5Wv0Zmtu/T+J2LWGPIRv4kyUJIiYpI2cXoUch13TwOgDsuy8pDRLeFV0
ThzyMdcmOxj9tk9NB0P27XRScCSLHgYjSTzmMW+GBDG3HbXzaF+YoyT92YDk2ILGoYH6kC4kpmEJ
BxUTVHkVTPc261yvXwmLto7ZQZMqIGwE7Uu6AWNeMUm4Zr0x04sFlPPy3AWN9ICnAuUpi652gTni
sQLrDYizhKBGUdjvSvZWdmnPvpX73YhI2m8yRNDEbHIeX7ZGgdu4zvdQSlgkKki7R9I0GqoADWIa
kI0IZE1PTsVAHynx8ntNxrEw0kKKOlHjbVODzptHQ1kMmzaSQtJfyC6o8NgQVi1DSZWMtZfxOwgJ
uIAudDGEFJAx6JNCGXOSVtGyMmbYkxcMvJw8rXWyrvXpQ88xOGhvLGnYN2MAQmkCqhwKy/37QU0i
UKf6l08bMfx/6948zlbu1LVEBdHwKnGz9y8bmPfq1fOMuVog9N8+jcuwFupe+PUe2pKTUlu9CEOX
JYwnTlDWAXAQo3h5MFAyHvxQI9lEXh91i7DzU79XjEFefhdDV5vN6qjKNJIGNckwQlYcMgbVVyNu
DsZB8I9/n1fD4QfwxFtttU63w6szgqX4rFoP3ec4XzzFl5Kh8dX6GD31H16s6LIn5AvtRIHRxeZf
UzAACx0EnLmr9FilJU4vZ8wME1yTqbeAH1hpFjURG0o8th18DylghMkcp82J6RkHtYx1ekoXZYxM
wYnJrNfyAm+CAVHJbfjMVGLfGTXqq/gubKRXj2vE1ZHGYdpU1tj724JS0TfJzDdGY3kqUB1/zCMq
lPgStUzy5vyzRGf5/aByISIXNwha65RMYJ4YOETQuQl6mIKMxSkxGGBo5CgfkKjsRu4YSAGiqYe2
Dsm3QTUneMtbBKXQkaPEwwu2Y7ysqEAmdPhAduiJbE5FvPtkKA+q98B0TTxqGvtJkemC5DALveVh
8KHWP/V+9UZe4ioV7W9U4+UNXmbSVYsT+EPqhNA3d6kqiO/xeFx1ABZYTGqTxjN3OPZuzK5q1vuR
BWhoid1n7IjrBXg5VR3TEgnOoO03BcSS4CNXZ6d+4DX5Re4LqWmWY3EkzC+rbZJIagUyDoqJe1Ir
bHbz9iTIA6/sNuS3dgYo7miTQCVSMcDTxiBcMHBJAcnRwhzcpp6QJwyZ2XHmHz6HN6PjGKjjqHyh
dBjVBto2UZxUp6u0ugyvmx2Ks8DaRkqZP2f/Fm690QZCpdBpYlNpZ5DaMMaou1KO4bX7GOv/X8T3
5TBFvx4zHzzFAvyM0ckWseE011dn02dTYyrhTRw/MnXnaIAXS5DgVJ/27xh9iTEKV0y4qd8oOjBg
dCIuQrr+pUrAlDApJX853S5cw72KkSg6IXbdi4D9B45rZW7SH8ijTvXjwGDlbIHVcaY8Las8LHQn
b7grvj7Xkfiiwh3d3O4GxrO6ivRJrv6fMjYrHhvF69O96bNBg3GCE5WZ1jvWoEGUjSgFiFcNlxbE
70QU9f0CSu/yFnw207f0m4H+ERHJCd4d/VXODiUlt2O5/L5F9bPLPyvA+uuKODbUPzq3VcEunYCh
Pnaj/qjj39CFPrCGn9ZyfVLPINZjAZct0+a34jb8Lv4tt03CPI11B7EsSAjy3jPwmZYVELW4rDOs
xGeumCPg4e5NaOtPgiqs5qbmpaGyqT301Xxuv6pAtFaXvh8XnmKjbWsxzKucnv6Qa3jDEqeQXhRD
Wkp/GPnFpQnaCNJwazHkMiDWdOnh5L8hvlyfLcbrderldwGYQSld1x3NEtjNbkv+3GFqqFdozOyY
AK9bUlC5X2boJzdcxOAspZrlOsq0JixxjHdMw2eMqlYt48NeBy+mcS5vvNyBne8xn/tKbbytW4eY
SLoI5+VpeW6+/KrQ+IMua1cCR8512o9+fY7lhFIhzzXsbb28pQwad890ZIgihK1nXfzzohG6CoCV
hwiEkDR8RlCzWKlabvjk2XCFRrYAPU3E06fE3FIOhX0F4if9eV2NuXwGmoTRQn3jT76OZUt6juXm
kZdLDngdzc508I/Db6Qmc2Rr3yH5Cl6aeSAOfvhgQ9QQxpXjoeRwXr8bg81KPqXKgZRdI5iihFZ0
YlaL0utnQFblLS1ACFE2lOK10YZoaeDevsskYogBZUi9v2EfbiJYT9WEqU7qXfwwjfkUwpgUYEDc
dm6rXYT45FT0YUBh43N3n2xrKxgbeN+tqvch94TwVqqsqRjz9iO2nlELKPPw4vad0g6+oaopan5R
BssypvN6JdO5d7LuEO6bMw4DzsvwQQtdqGzRp1cA/JmUWZyf3LiVz5aNh9uzn070Qwt7MpMZ4TM9
pQvei6En+rurLv8ns7pS1lHGJL+FNyOTOegEOwaddETF0KLjmJrbz2V8RY7adSLpItqhJcCDCzvE
On57VDXedk+zQvTMG+RULUpUk5mPYE1YQ9cwZz/9R9Jkd5+cpvH+RA/iV5UfJpFoFvlQNsuIquuh
m/oLWqCUutISaHCsUP7t3WyDlLsZ9QYVW4GO5Sy477Xk6SpqUXQccJK+jx5XLLentZVQgc82NrhA
5K7r+wF+XLNfHw0S0TsqBEiw9jpR338FslAaRtpz6MCuWJzg8KUGN2L6xlyJym+9EgeOFrgG04hS
368IvQTHACXQhQl/yC74VgK2Zn03TCtjRix0eaxIL4o3LanPurhTO/sUf/BlcrKB06ptOehYjuPU
lizkq5YSH2T0YkcSTsQpA5OGteXPgIyiyWzTFf1BU825Oyah2R5OJWuYL8hTpmeh5Cxm7nak4rip
6fdo+cFZbcv0v4KLBpeuYCds8GxdCwQeieKDs+9pKYkliWARyvpiTeNfl4eiFd5zl2jlIL3MPSHb
MtpfjGFB2L5scccUbHytke6tTpDOEwTF+f1kpP7TJBkbidfGx/Hg3IfetTDkGevrZpAsVG+Nun6x
ejonBWncZOkMgxkXMAxS2j+O8iGBavQidzglta/Ull3MiLXSPZRc6Xeq7v8qCGREKaf1/O5pPf1G
/8yt4O3eavfv6F/Fvuf5rsL+lWSaGZajcbPlYWEZ0QxFUyTXVnTpfjO7VvX6yshPkUrGCV9+BaD3
2UJ8gVrOy/hCHwzkQM4DUNpxTa5AqLbPkOm0ogBTb5tTkRIszwC0gDqxiOcZRk8RWE27zo65GcWA
09hjsmreIncm9+cZbhbBLHf6/rkoqRlCObXXCd/uuIk+vmXuuHkd3uGVQyobDgsSt7L0KNdHm/dP
QMND+k0COj2g0VpIYlXzRNcWmPYpyUN7UNIhOO6yNnw1+ijuLLaO2vXeuhdL6J2KrOuUgrX+1gRH
CELOMFh54NoVrpvG+QJGk9uu82rLa9cwDKfD8a6h1DjLbg70qZitRPYp09pN5hj/M6HoE2PRzeHL
lTsMxVVUZSU/OcIOK6Vcfr6Jr0Sh0wa9CaQYX3/R9kTTHkOx4+vCQ6l2+SV6DDPNNXk44W33fHO1
kDZy0hxr9uhZBSpGPtsq1bH5gjnC9kMMP5BjOP/Cs+2vDpY3HEK3+AU6nz8ZbODzmetm+1jWyYZ7
z/fY/T77/7je+Gmm6pVkMGCjKcvpUOWaduADA0n0tET9mCFT5lFBzleXpZPa4LkmTCOx93Vfmxkt
PMgCP8Ac+fPeciOIiL4AjeAI+N8OZMIGi3t9O3ZQ2DzXT6o/grkqcTC/vKUgOhCVsKl6ftiQ0iLG
odxY6Kp3m229uVaG35CQ/oe0/3l9cOLiu/Oaa97QAQtAdGou1E02JhQsZ3dgeIXjoWu+xsEfOqZc
YVlELG1iBAcgViEdwKWfMF3HBLHjUNEfdZ7PwFU7o1fkNSwJ/dlVYC6+G7bqzEzdKbZZLZyzS1HF
pGgaiLNMNXTflFGQe3oyyyIe4gywXariId5kWLac01BxP00bmGDeoMQ4vDp3qZnwW7znRPV4e4Mr
nGWWpWWQMFBEfMf+68tO5Zp+HGyyPm8W22QzMe/CzQKaAx+/lcb0ncFL7wOlgkH4KHwkayBS8aP8
QxaI3fTaqPXz6tatuWK+LszICgfOig0ZHnFBZ0BsjPVHyR9iCtM+U1QMymEM5RucA0cBW5D5bX0p
dbmsYuhBpZIydIADAU1Z/UuKhsPAadCRMU0+b2OBxD9cx2BhZ/800hjE2w65lW7t+fln2/0mu6B4
HoBZme9OnGH1aWa6bV5Y/zM/5GFHLat7bgxC65iU5WdoxIVlUXonKREyoKKywK3a1D2Oe3GTrbqX
4edbxAddx60OTtM+A5yRAniSgQ80lscTjBL5hdoaR7s0sdTLFliL2t1BlhBl8SYRUGv9vg4aqeuZ
PPssnqjYHIHiPKNu3VReVtjapxHTrYb6nZPB9D8BJW8YecbureH2SJgS917gyhnX+PJuMkE0FqJO
AueZrvMrDvfMcnDO5hUq5d/x12twJSdKscC4rM/NOC6t7ZYmFAP6q8JUsghk5e5dMmRnHhvKfBF8
XRvZMyncBN7p61OLrYrDdaWnfqYSxP0tRIz+osZBgAfOv1k3ihaZNDtt87UdPu5Zo3cC1fsQhjkF
dhKGMfhJfVXqm3ThslAqQJUNM8bTNG1/FPjByYun2l+KWd+kWaLVzN5eO4kWkiPhVuF+b24iZ4J4
8qBRAOpaTHtF8T0v8Ey8oOaJpij69ivv1HfVC2BT7UfTMLXCf8adMXgb8o1BYaIKH7jX94d4iPeR
Vne1BXzQv1SoG/ztm5jp0jN9cunfUxg8KaoRDg2ui4uaJnBUoQjZNbfXWAcJ7xixJRI6WYNqtecP
RLpKGgLWRRQN/ppVLouBztSDVGyVlsQYK2EIK+6+zSC0Zob64suvlzKZxg5yy/IQddDsx/TmAOM/
O6TGn/d+1U3JJRHVf14iElOMh7+a6oVTh4DoNSCy/oysfNyx3uRpfjfKuntRimIK9+Vl5L0VGWZ2
+VL2U1ZQ0Tzok1KKv/pOVjPRiIYaX++wHNWiAX8C2idV/kC8uf1UHCYVxK03PgDahkp+u+3NamHS
QlTPAhSlcA7Q6AfoOIdS7w/lyj6z7bF4jwyK45GlAQiUaTJh6anOijI6+v4YXV/t9+4eHAIzeYKC
xerP4pHd1X6Gjogo82RE22eEr4iC360egF5Gjn9R/nE73BE9Vsg54RvDLF62FmTxonoJu+dKMNn5
9GgirNHVGcKjH9XrF9Iiq3nBdG+FsjOsX1knOarUQY8LYct0TdM2gU+ruj9pkgvWqcyoSjdO5bUz
MC5S7n1zQAzEY9yDBJpnMlh6Rj52mx61jdR+wfN06ldMH283Aqg6vkw8nU0zK0YoKTprV7ckXtAY
GdnE2AvZl9ztJdHH385rAROCuXfe2oDKo9LfSEV/uV5fvS90OQQjHkUXtyC6wSeZzigVAtiL2NmT
S91LRuOREdtWmtFSv+ZwZJrva92uwXrwYYtSi47QALwmk9SRzBVfRsV2rDSwJvqQ5NepfWd3JJRy
bqTXCYAtF/r1A9NOEIrnc8PXySFqEg/ULLD9D8+XegKB1CEAzTZ+5mGUSAnyUL557i/1tu8PyXS/
6rN8E4LBZCXac1DGLlzyvgelPYWe5aXHEZLVFRDQprgrVu7PiCaslMMrB6Fk9uUFww69Z25nOtsp
Fw16XcAKim87QuLdGZW7Lpul6p5DFMJ4ZA0hRnqZdbVaBtLTHsHfozc8OT5aDKUo7fGpms/lVtpt
seIIK0O2QCjz8Gq9GJrumnKpyMXGVWwuNwhllTLhzX0qYIxiG9pS5MIyxEE8R/dRdvfAs8ZIRF41
XPWwYlTIpFHWzIlVGDK0zmMItJGoyId8bpZE6qUlpuQwgtc7qWCGS9DlLP55X5+QZ3anukdI3UuS
eoVrDSYKJsxYZTpi/bLIFnA3dVpvawfb8IHa2brc72zbsom5rmyHaiMV03yNpCuR/bQc7fiLo8fa
stlWAnxMrhznyi2+wHhIPIXC9O1cTTk4PWRC9hft3Y41zNyacsKtxhAXoqOlcIjpVKPdGrQR7fmJ
KIpQ9mgTcgNmR8nLE7IzeVwXB21se62xrkiPC1vKkJqif3Rf/XryxiyiKuX2utMNeX+rbY0s58pR
Pm6bAm7zhwvdHv4ge+zxmstNHyU5iKSWbMJv2O2K/LvytseE4Jp8Y/2B+yoUbjSiGRLutTqQaEST
ghQnGOzEBceEbHgz8bpu/sSvK4LVUUQd6cVIH8Gcg5xON1+Xw2SKgo41x3KoWyBeFqYJC7Zizajh
RuLROZfWFtaWCmz2kBz3WDTs6wtsqDYdmUGtQSO+zBBkx0G/yxZK/Bp9VSsxV6eVcc12fM+z1dir
9Latw4FirNmaIlJj1LsVyCo1Af42/QcoEQWlUIfAFewMNieV9mKvDV79iW8LtaRdOeceQBMvom3C
xe2mRAFoq7w1PUN/Phi6fL1DnonDN9FmJpq79vAxqFCsSqW09I80VZjUjc919jpDCf1XZWtbGkqZ
pIQ3R6RhZbl/N0bw2xxcGvns7KtjC0kgzYy4o0VMkVgy2zW8r8LuA5YnrPw57nZs+z25M+J9E0EN
tcd8queSFFi3f0RWsediQYXyyCij7tKuy6cSE3f1BTjjrrUYkF/05Geab1oYzuGeTgDihMHglxxL
bzwt5x1EuJq5NxCr+XdJ0NyIQTK2IdIL7v2pwzfa805YsUbH0V7CkwHoM+ly1KdR+fNsvR7AdSRn
XhDaDZv/J5+/eQ5jxJi+EYyadlPhYQ0M2I8GetBRmG6zIbm7OTvzD806U+Opid/6VGTJa4JDc5XI
MxdRVkIxGKju/aIbH0xJWT9imoai0t1djuiNWLxtlj7r/J6KY/H9tDwqU0P3yysxE+j4/VXV/p2o
9T91I2ofaqIbHWIFbZrmMZbMSet8RPTAymm7UQ1ec4SVwfuY2VhrfG4UZjlniP1ujDeGBpzmf27E
t0WCEyBrKuSuS02rp1R0ywilAXoVWm1aDvTIiXMygJgCXZABRbwSy6Owv90dVEklDXfPuSRqm/YA
lL71x9nSLREaJg7yX8InoPHRRySEQ4CbyY/33+esbwR8CXlWgpYZq8jbbKcmEMzSBIFzkH3f2gtV
CjqoXtDix5ROcn6ooSo/DOiZmJwf+KPtHJNzQlRzeEsQjjIL87DXayEzTlrLdArNGQeRsS1M88qW
ZT1XKGHiX6EPqzRJ9SmT0EVIuVtMvxCbKY4ZKKgot5ZVjhH2g9O7HmsWSs8afIxCcUlx3zWMiXHw
UuZ/jzNiCwnROEsGl/uFBaVfS3NflBtzuqbz/c0KdwqVESDjRj0+IfYkW5BRUlsQN5LSSvqrV0lL
moVmqJcgxiWOjprajEbY8k11/BpgSFzWPDFEO5MVRyNGArdqedoiEO8xIJnFwdPptQh+puktZGOZ
H63Ef8A26lf+eBonGbB21yhsXEu0B6RPvzhjhGCAwtNUyTNEMF0+PENUonWrFnG6/H6oDmTBThIR
hpKRlVcA6BgoaDXeKKGVFdKcw9gNIYgFBvPUm9PrZ96SIZDDtYVNEgWWMDyfSHxv5axzj1YxExOf
fV0/Mm4QqNzrFftsbZdfZf4tcWMVEECmHJRDLg2mhSc6hGbAHl2p0PeRLhC4s6zp/t2yVqpN3u2t
06Q10JpNRcvujUhbsJ0aq6QSV4ZMiYiffkMlpvqyAEMfhcsIG4K/BZcJmMHlDiO0cS5D1Ggj6kbB
egAiG4eDuIcHwB2BK/6AQcHKjm4wnkn/Bd5GFGY+o8q8o4LbBZ+yXY5hHps1bHQ09RxwPQUrvhr8
6gRfaqrBao5RoHCxYYVjcLuDbuiFtg4HotnOr2hBjZRRYjVeOcLbRqd6bgMlIFzcRO5dXf43Ripv
tGMQ3ELd2bqOMb2UYpkwEmQywQX2Com+8ihfKOCEGqAgb/82SD4Wgk6g52nCcGo54FvzKHdTRnMB
MeMGERNDdcZ95S0ZNcK4/6MvVGqLAxbtyXeDnu/f22vIP8oE0FWtRGCxH9/4/Soa57pJmClI0Kj9
01qZEX5w34qk5rldA9qtSeTPAbBugNVC8yqFCwWUlkhLlUvXdmV6/QeOjHFr+rNOT/3Di5mpB/5U
5GUHZC0U59fh4v/eRytvc70H9oIpCHi2t+bFQgPj+bS5hR3YrjTJunMOd3ka+L6CN3SEYSnAD3oU
76i+QdlKCSE3skbgS4nMgLrZ8+jvyMna8Pxh7XT+MNQYVB9Mxq+BlRC1cJXU7HtqbrXC5uSkJETN
c+/TwZMIzoihCW3y6PhaebhZZ7MOwg7Qmz7kDPJdXb4mcoiZdwzkS4uyJc0zG7qasZ1XeErllfX8
ZXNWiLxbk2RvBECHiqJmmPkFNnTp8kkc6EL0TRSodd7Q32IyGMIH1hxVcihqqWBy/kvtYkD5396x
Q1S/zdf6dZw1pqUfD61/cFKI//fGkqkPol7cNTE659f10gE4QsAF9lZPR4OLkK+lL1Wb8esjMtnR
R3FkNKBsNKAISuKnazeWo1COhjhwkCxv3y+O1RYSZg3PXEu9kUeORqBAnXATEEgcbVsOmYg3V4y/
Docu4GitoLt/H2qwCqoxeXy5QygviP/IPXTmBkS6JZiF48Lcdz+DY9bhvyb4fl9bBdbaoqo/yqJf
SZvPXXhaweJ3Tz2nidwX8moMKKbdIfBwwlKaHzAM52LaLl1JYKB+ldjMeAKGBFuqcae7uLw5VcGZ
c949iUwhW1NgYaMLcKEU1ZXZ4XND2t0MtflIB/Oof9MHzFWHsVMOpEMYCPjjc+TiJEZU8i3S/in2
G92vBbq+fvilaF76yCRlUnvEbO/r839UkT5HhpxVh2KqsBpshLVCJM3v5TEK7sBQ/4WsFBJPngbw
0EQhPvpkbbkCp0Un1eFuyer1ysb1SRLY7ufw5dPV44no2fIyLTmBl50K1+MUg134Ix9jF9U/nZoT
koPERx/hm9S2u02xZ+q6vLBLgW91zPPpO35FYn3SywoPzxRhNEdjmnKyFam0IjmULo2BgC4NRV78
fLGIEK6Gtcwj+yuWoXZ5PtE70lOl2sMjw+Kue/eu51Epr+qc9LoGiKMsBVEA8WrCdYyjGoOlC2uD
WuZ7YJcLjGuFKldyfDXAXoHdkaWqddbTHkV2iEC4w3H92g4JzocpB5dse9Tp496+Mfr1VGo0R/4Q
2AxCiB5W5IiT2ClU5Mg8WkH2ZGKXbbUOXfW/ORg/zWxHodeBqxIcfGCCalxJtt8rnHN3PVs8ApUq
COVQdxnJNKgzmgn9gqQ25rxjiDrddTttXK9P8cpjCBKp5SQZpg2MLH85tZqB57+dD8zTH1gNc9Zs
OMs0bS2enMi5m5rOFf0VfNRGGgjTkVfBNTpDI6DbGst9jV6IcwnC4aNfBj7l2GZ8zFMI8MMJb9Kf
kI4QDBLkApaNZxD60B1EXns13iisSTRfGOXNR1dnU4JEsE8lYSrmRUohyjeDVfgM1w4lyZegJE0b
G3knaQ2n2QOR88CvA4hOLzJMJ0DjFA4WABT1FBCEZDsk5yakiwxODHsjRos0Vk/5uAl5GmVoLdvz
4c1Q4NxKZrbEoPIspIqteFUYujlBm6U2HnvZ7D1L022qammOk8jijidfzHkbGuDN3a2I9SZWxjHX
IQCDsbW2fMPFmqCv6o/8Qf67sXWaxek2Htif0ndVt5j6A63WhQXoH5NOv90X8HIDFa0VSODdVNtD
btYjNrxweVoMeZC2tAoB+rn+utqnu/rW8RPN+ynZL4lk7Er6o/byb83kGNcYG5OkvfBPTy62o9dZ
LTGbjyXsZ0pA43uftpdPYLZzn3P2vvUvTBB29I99ajBs+QNZuMdSX4LWmvGcXlaqBjbBZe1KCHIt
+ksTlcnvrr/W2le2Te+wwQAD1ZCppw/YGv6HOFSBZeo8VLR3VX+bkm+QU1PHLDCKJ26cu/54doYY
+oevV+b9m3DxmhtyWEUF8Sk8s6uztHGMV7M/zkR0kDOcPCsOhqbx0gwJSDFfoyph+ym+54TMAple
hOZKhC42ZWJuktHpAgBeMwLaMrCdJ53Y217Gw8C/gSZ2XzJvVAq1BXySYRtZ3TnJi2sT/6tER2XJ
vIw5DSQraYuUqdknbBsJQGXxeLgNbYkHQjMgraAm8Lc1oWQOMgmxWLqymsa71deTouB6gCOzQ6SG
7tfA0t7b/e22i+1ZAla8X7svHxPxueHrCd+IhUGGZl3TfrzbCTLcuqT6u4scBHMYm6kD7AxaaT5R
gYecoOIOSf6I209AsUTRwsAMgngkUl01d/8zpbjhL2iLo1GCPu5zRGosG1OcqzES575gjrnNyYQE
OBys7eM+vWkyCqO/QEtuJ8Lr22BcbnB+xPOUcptcgVGQH/bvmlb6zk1mC0t/D3cbqgh8TD24lIBN
D1qOzVf0mF6Y2Eo3jQalfhqqIzUrzDKEfshEqWPsfvxPescyY+U/57L3BCQhJEgy4VBC/rDjt0EE
h9mIbLGuPHrpjYnUQpdnRT8yTTRAmEAKWxJGz5p/Wog2M0WwI8qqXjNvp/jTC5fkamQBDkhZub7R
6fZSrH8RCeU+LV2JnQyUm7wWrfKoYII1q7G0RUagpFjDiUA7DcEzTnWb6vENGSWPD0zPntMWkAxX
ZmHbNiOUMNN/rVQBpH9DFLXURj/jYpPaVF51S0nyC2nkTYuXSVGGlbELN9o5ZN3PIQbADfFyn+qQ
po4AD+dJwOCQ5ThHYKn+UQN37GBgU/B5SsPkDopVi+aAgYAAn7Jxu6MSqd4jzep0fGbs3XMo4LAg
7637b+RY5GMgdgvn99P6z4Z+K5JbY9njLxEZw0yi2j1LxkexBmXihm8LjTb4n8N1c42n6bKkpcj9
QmF4D5IxQtZ4xslbP2W3ko3RJQYlgx+ITzkPFpcaF/3LpgdISN2FdoogEML4A9LLp/458OWViKU8
OiYV8rPscbiWyX7uyvKI8cojIsMWnhDJjn3yKSfK+1KCxGE8WvTWyaln0vEgHw/HZj/Pyscj07I0
Kw9sApiNV9zxEF2R5kKZRm7gdPpOa3kteXzVkQtOgYV23g3j5KU3rtOPCtCQcJ8Yon/XQdLpQN2S
qWuE3CfyS+Fpep+g9MRXplEIE9vKd4T6aGRv6Ke/Yx+KwpXC9cJTkksJNhaRuvWxVY7qKhPIeq2K
V97QKVYHg/DT+zVE+0OJe4Tjrhn4Wv/fApUy23wmV/J6u62+4MUYdBGz2WnwQv6IL0yNwQITh0oF
+2vFuVirqgRTLAwu54YKYZ7tDvKOJcyFZyAypIu4/y3E1wfSAet+5ipo9Tu1PsrkyHU02L6sk/wa
w6cxS22NwDSf6094pLCroUf64TO9/YbTGNzF3l7DVjIfL9PKUnmjG9frsu0IqXdVc9hCSiEqrS+M
Vw0CF6XyCZHBmqx/UWRguPsqwQwc9dsDIDytaTce2Bkn5oFX02VmAauCm0C7ne8bZQmny9L2VSdY
wRzvIS1wFfYQgjHDThS7iLbE5noBuehZQ9JTBRS+YrQAUYcplwh1ygPsZa76cTY58cZtyRbt9woU
upZk1LUxa+RJF9cMuGEwEHQ/PF+vRFzcI8dUxMeEFTeJJKC/xhrU8m4r7tKyLelc6NCWoCmDN83P
3m/2T7VdLiRhSy9aCu13RbfjR0aCrym3UqQRABa+5pRGdwcXTnq9Qg55RXFVuuNCj4iNjXOKgBbp
dpS5NKNBIpNGO78yAXieOJ1w1v6TXYqHXvSZHVVY5IAMHeM1vw/OOVRhqfBR6Wo6RSZQdhX4w99j
TJcZE/GlkfM8BrNkl35wSwzg5ibCwzh6O6B+U5UjVC5IqLKzifxP74UK0dM0pcBvQxatZmLcprzT
Uf7qH5ZtZnWpXyi0+3aRr+SCwnl8CZ3+CgBC/AXWAXnuHDviAHWZJv3pZgsICFmd7cqtrZyz63v9
BowgOlaIaaFeRlE+e6w5p8wja6GFdgQVPAfSfw4bU0vJyyh56ELVguK4z5PjQjjSeRQvBOHPmdfK
K1XKqJgKYSXv2VpmQIO444LoUeZbhUcG14/axJC1NxgFDQdPkW51UVmj/CJH2eLtxU8v2flb8riK
a47uaLo5DmJy2c4EETr/4aeOpsUuVztuzWudAtl3sbjzPyli51e97tbOzF0nw43vW0+FAG4TOeel
lcdhR7dJluadJ7qoGeujHi+tbB244P+eEZQiKPjr7YhAYSlIPMN4T/zdVYiRH//TBqEx8eRSzNzJ
9nGBp0486IFZnrAENBbmAoeEUI4djGqxDQqPE8eKPFiGSmYVMMx3cXYy8AaGt+V5PVV9oeQ8PCqv
z71ZZDkSf7q0AO6q0auz5VoSDprxpjZK8ppsUZSJaF08WrazVAnvz36sesPkEGUrroCcs2W0PpAe
8U1Iw9Mm5YyA0fnCDxocchsNMPBHX1G4XrSEludi3SGB9teg4UchCZ5KwWihC+mWjWt2/LdlueNl
K0Pol1/bvFT8ULajWRdAlE73hh3iE3M0jjpdqPwLnwLxlch/0tkra/Gs6MzP6+MvmiIiyCQjrUPE
WVqMfocRw4lna9N4zuv+khHD+ztKE3iYXapFvOtH8k/xxIFD/Grya2NMzCsdHBEue2VRUiWEYrUI
qsmTGC2iH0kpzdQ/5tOj9Te0kD3ZEXBr1Os/TPFF4vXUifu3+I38PBOpQ9HX9losdak0HRXA70ra
ndnwRCwogj6NIy1TeFod0EN6dfNVE1SkFHT7vPsEt76pGXsG/g6+dOEiQbFH3VOjb4G+O67mhxBe
rg7f2DxsrxJuAoAqJqDB76A1TcsC1rgFlFKO1dH5K5JD3JMxElW+fzv9tzrSNm0manKASxv/l9SG
zrj863Puhl+0p2JeRXvrp+rLIN0Ot/2IMqm4mogqTToZU/MScrUwx02w4b4AF6XIcPBm0gKZUloZ
fqO49L3AQ1rrwgLuEKBxtp1jmmW9bpPVo5yCg1PvG0drSc55zTiNR+hwccE0CpCR2TNVaKmamLZD
mW62gp1gwEc5bzJcLSPo8//WnjuFyyVsmH7TFcFsKypo1l419ICw6p94/mXbcGF/OO8c8YcSsaJx
9wpfo84yjEozhBBIncS5iXB7HRsZ/sxdJrTX/8TQ7PopBwmmDWmoNZFdENE5y7VPwLFckKsk+U90
dZXS6FiMP/TNIPOMDPJYFKUU2Aks3eBqC+p0kFnYMYSeLMvBwDtD+OzWWs82h2g6TYiyiFxX/43b
XgPWq4fBfZJuga3kZZxoPJp3Y53M5ZPsCuKGHHLizKULLXBsMi9UgO0kZM/phCKz+HZjn4yC3ufS
lEQn/e58R27h+AcvykMBZJ5KGHCvqbtZWsv1bkzcG8+eB262ZGyML6MXW9hvRkrwHZ3ewCzKbk6V
zgUNGeiEZBx9S/hZyUmYpmRgaUhbKZLecH6hJl3bOzJD2qr9OVNNI+TsBXD3BHtXRiDByGnagMmE
60t6I2W7VXHFxjOl1WqPWc58I3mjshKD53Fd40idr8yUEOaO+vwcxupF2GZqAe6/sn/mRFrJkI/5
4yV7HDY0TUO9+hiLNfRCioQv9UajcUOJeMAH90/tqtjeK/KfhhTjy/erYXO81Qnp9TmH46SuJk7j
wfCuRNXmAbvfdjKB4xavTKjBmI0UzfYkrutbgNGEUR1ty9PbZzzO+1KqRg9CHvcyIddSYlPvhMtb
OVIjx3gIWu3sfYqJG+2S4pKt74DdtAexhh4CbR+/yfDbUJrQ88eLOtfCIi5lj8ykXMwIfMqVHMQ3
WFBk+tNoWfMdPofPEi4SNVsYtEUvtkUeVdSVS/uoUNYl5J/JtKJixrwDzMM6LMwnl5EqVTxxUf/E
j1AjnfQ/PhJ+0vMR17Z6mCNzf0h11zLmw/ekUi4aYSn7rU+BefEDpU45D6UZ3cMwvQo/NBgt+Bs6
GCg1Pv/vaxozxOB9c9cUhbxbluWf12EiyEnXkUDf+jurbHPixfs+XldYXLuCJ2pR81d9BXNFkmG5
GZzAsYkBnOftYuVxca1f7B5NrzLTmoM2VnXMcZ3gNtwX4yXlEGywK9IFvE78Vly3mxRlu6sk33/K
rYbj0IPdGn0yRjKsQ8ldPLdbIe9XPtkLYdqFYLVGqRGcJVdnfj0pPsHuLH2tHPCWcORciTTqUvoM
fiu+t3iE/Nfsu0Ly6nhv3vRTkAMzxUK+F8u4dC4mcBfpJGhzOSn4ft8/ec/v8fu1gj3oLmjrXZGu
sJ57tNg7kY0PtNWlLEs812AsHLQ30xbcLo6SwlJ/P/BdEHMJWJyinZEptJPFXZDc1SPwmHUtoQwu
YHqvQM+e6rH99AmJ/OHZPkRU0J8eMF+U5hXbmacMpKY6Yztk9MVviZV0gdqdqOA9lxhvqddaSAZY
vOdjNM1UVI5LNWw2vcihWzDPOW5DDypq/znj0AQftfXvEOYN6ukMKvCL/pvYBaNfA6jjoQgGGtfo
ETM/gDn6hKYQkD1EcAmcpcU4++NU+sc6J1ZUyVPmh+bIvC/7aGcTCM1ac7jAEkycXVw9J+g9ozmK
iPkSgt8V6dMOADn+y7X0tAHlae+6vnZH3/GQfv0ohS5uogSs72Elq1u+aFxw+UJiHDdlYkwaMt03
irkPd53QMDA0Q7XZ0ZJNbitx9xWo46LPdROIql6aZxbVRAVOMyU8GOPEBDHY2+uWg0aFwWGtVrGP
0WhQp9+cu1M/0kv0V9c7In0hQ7OochO1SfcGc5yc7roLVJOdrhfyAiMV9prWT+2HvLn024GDpKOw
gPQ8yhfBxX5USRR7GlHuxq1bV0r2crz5SA4zANsm+LLPj/bzkJ7jJNAiqkdQXY0AovNousURDr04
30mqPcH09Nm/4KGhySPwrV92ct4NIosNY92HTqm2xHsVCeqKrgJmGq/9Pa0Feqav/ir2eUaAEkgH
GFe/iVh9/VeWCyiFJEZkl1Cv9bK3Zame9Ldg1XgXmcgnRQ4N47m/GSQmajN6KygMlziEWrokTvLF
wchEzxIYdLj64OwaeVqZoBYdGXS5GcN4arwoNZYJizsBFNavuTPObHasFFh+N9s2RUZuPCwKmnL3
lhNmzgL5JCVxwaKA7UGcnsKtpkh2t1CjypRgAmBPD+3xZuadkAewqgRpmdnZdsQRT+9B6fTvo8wg
vxeZBOjEyfS4qTfy2S1JA3PY/JJfFgdHe2nIVzzO40h/MUp/ZV+DKhSpBNUjAEWtewx/vkZZdP+z
D5Q+ApJpH4FowA18Sptxhg+p8ujljSJfNszDvmnV0if2/kblheK131xZI6Ntau7I1hCkmhFvfGsm
8yGNARrbkOp/dWD6vOO8sJzMeQzd8USZPPdj003qlLENQAg3/yr+skjKfr6gRVSvzi7/MMpt9PyR
MrWafE69tp2RYbP9hGWc2YK69P8cEKt2e+ECBhwHeqySuCwIU6rMT1ws9+jhoxVN4ZH2v1o0tAfq
RPhToF0hAtESlH2c8F2yLnDud9Mi9mUtNtvNHiipPA+cVZDP/SHs4MNmL81iatb+r+pHggjVOF3X
bnkC3aUVEhwy1+vrS1xmpSz3MhocThl+LbUA4yvucJBr29NROLi9rh75JJ6lfdDFtseO5BujnmWk
loVeQQGni5MkR/zuKPMSGqaCN/9Svo/u1lhohO42xcy7NMg+UW3MNpjKXb7M6a5NpLOS5adRVv1d
Lj29NHiz62fnXwbzuH8TTKRueKnL7Krak7I3S8KhlZokBjHY2KZmuPb1uhh0dpbR8AUom0teGZvJ
3eVIMoM4/vszYCXvqRJWyFK042tILdtoyIYNuZa6qYnxduw+oruAGC1CgK6n+zdmFxX8qrrrhaFn
zLpg6vXMyft0lizr2lcPQfXJl0N5us9iM1ek9yvxUbwPre5vkfYP0oQfn4g1eZ7bSbmKX0soukab
gqED5OXooTGbXW+xgD6u/ac8yTFN3TSXY48JTncNLw++rmsH1rwIrzAYF5gnJSvfRDtBENRplICX
UyMdk7BDQOSCog9iSUjlv0kxBj+nhb5TktOXuR3gIp5Nqfr/sqVEcoaics6vmw/EJ4jhebN/Am38
Np6gZMw9r7ADifRDXsIz9hkQ/1xVL+atEceL3/kLlRpHjmqHlNk+Zrk7PhIwJp/7yWFo+qOsuQIu
I8XA+3jdM/ZgmpPncbM1S14Jmb2ayzG75db3+o9pua1dyRDS9myJM10SW+AO+ptQUDhEkmyDOxwm
x2/g6Fto8vrOHz10WKI1FZIVh5z3maijGP4sfL74StR43pVfF84fKl+t/EzEcYCD1SWSeUfXyAmg
44yy+k0c8ZsO3lJmf8trUsKfieL/dAIQ3re29GXneczh0uPjCbaD4C9pSIZ/2s1fGZ4RwhH0h0GW
ltMewqZ9pPogOiYsu3rfQR/CkHjlcQTZaG5UA2u+84keiQU20O0BGnTlLW0hVV+2X9JtsVC+2CI5
K8Bj2b2h0Vwr/zLPW7/hX2iK5G2ceTgEJVKqfyp8brmoO7JZFImHxpyWfmZMp7nYM0XMiEdTvoHD
m5GNWGOtLqSQFn2yj+NLzJ2LnL3HiuRiiv6rh560cGefmQyyV9NmdtJhtNNRDmembebwSOCTAtyk
QLjulNuTsjyL3EP5htf+qJADAFpWnqaqlT6fDktGaOcPhug7EHmcHWRQakgJHiigFxfZpc6kcTuv
VwO3FQuG2x3i9xbxwU44CE2k1m5wjp0+TXoAYWWiLgddufysiu5fh+fBCBOsTgmXDa49Ttg8o7Y/
oOZP28nmtArkbBhLMZ217CuOzpG2JPHvPigrJfe7YMCMpW/yJaLTdTWErFM7wo5ioZj7DadUd1h+
LkFht6utPYTiLy5lzLqIZLy15q7DFVN3XFPhGMFg4orvY1RT/lhSI45h8pRIRrHsQ5SP6gPJZEsE
X/dBmk3Aydx4hbFvXnyyWIZuLUIrUEPbX4xzppwToN/2VDTWw1jma1I+OYbRbaUzl+nupgxNhiWs
Z98pO9PPUctGSSTUGTU4I0cQIeueZd/GL7cQ4Ygf4wUnc8VRJ3C6MZyU4SwoN9mfUdW73kdNvP4X
mPnVKFJJdWakGFJkpWs52r8qNJECU8zjyeXBbyBS0ENKCy6QVDutu8DmKNfqzQSn2lEfaJEyfMzL
mK0BckrY4KjI8b6bYu25GsH8khN0LkFwWLEJPlQGwmN0Cx4Md1Syj43Ce0ox73wjP2lXoGNcaQ5J
s6zwVUwSkaZtUtx9HTQbQTOyJblz2+rwt6wZfP3if0WVD3hhb0BQi2T1Lb69GFN1MOTReLp/7kFu
THJX+36/M3A0DN7GKMTA2IlUXqIraf+l4shz42JqbShcKkw/WKX1Wu9LGfJ34GPyNp6P7Ty9bp93
D40sJ79jzQTOv35Qi+8q48sf8IH/8p0oL7vEDniZLcxmZSvX2BX+5hw1uxnjyQfdaqaufg0e9vJc
/hAxrUBSpnm2mqA3qz7rJy9fLc+25ofPMxJq9+Y2TJAStTZJOKJkWmX73EyCV1Qq+GzxgzyN0tbi
xBpAzs5j+2LWolzV4ramEOxTQ7HfQRw905i8YDPbrDklr1FlDMHVis0ZX8j8a7hFB/igYO7I9jJU
mfiNEs0yUiembhWSgaX+UtG7b8atmtoMMJ3pnBQDC3PHYEs7TknQKXDAW/KpZzr7QDcVe5PUFIY8
0FPjgATKoRz22H9TJpCY6aXsAdgmPoLt59v8k2RDHDYU9IPRU5xuKux6b0GYTR2S9tCTkbwmd9xa
JK663zsgqeyN5OSGNikJ1pSIHf/0YemPaidZRBOmzPy/5bWUU7oWPQMvw+NsTJVPGZy/4OCoSHYN
gGXC6wkQxbV7mXU7X5znhFrlZChZdeknH706y4/jeQWgRHEBo4ljNxRCszrmkzsY0m/GRPUhRbo+
nJD1wuRsjPK5t7T+9nYGtBFDKh/VU6IF4Nbe79Ys8ktWWIRnnO9IV7A2hzFQEjDNGQ9/2V3tmVLB
MdvSlYGO6N2XkZbxWiHFiQ6h6jEmlJ2Rtvhk0lBkfXBn+DiDpXieYwfxB1oip+mv2whi/RkGPmbB
iwzubXRT2btcehDCyWHhHVRqks71hM/zDwB37oAQPpTVRQ7tA6E08mIMPLugqyKGkgRmdh1QeH+P
2tzZhwVCcABLIqUFNzYwKYCt8kg0zPAGyVvEXykPY3qd5GSMDsjS5wU5D5mMdgqiyt8V70w1SyEb
7afV6NAfyJGF611U1BH34D/L2B0iZ7vRyEf0d7oQJ9TluahvJhwc8MufP1oXiu1nTVhyKs923BkI
fgeeSvM8VS61URJ4tbKJfjrx8WX8d9tB9Mfa01Cw3PgTpmMS1si/0qSTpXDX7o3VbqNABl0y6cdu
mRvgHsQNL4QJ+66Nai+JP/MPkq6V1PMI6kyWRj2b1rAsohcSRTHXQpS8PbH/cb8gPWnqiHdLFWE0
L0D1Sc07Iv5uUDRV8M6qmo+WNvksrkO5KC5Uie5BCKKZOfowwXDK0KxERkW+Jq2amwH94X++80mX
fBTuk3wY6BlC8rxJ5jMGoJy2/kcCwvGujMNRdretzu+BZiKFWhMO2Dgijz7vf27V0Umy7HH4COmX
h3v1ZdgKgcTVS7j+e1t7alz/Bn2+MilS8eB32V76nhRTP7e/tanllsVZRmbvn4fokzIhf7n3IBvH
GCehEPwIF1eOjKNaXibDeYo3El7FS+AdkvWf6hvUWGbvnonW1+oLbwGlvjs5MuH4oSz8tiqlGpWn
s83O236d20BwseDCsuJ7p+CRyhCkHEnaQHQ0kQ17AgjH4D8x+Hf+7IFGJ48H8alOkCslq7oL0lvD
cGyGMq20M/BDZ1qr6thJHef0lWXgG0xvVCuLNj02t60fG5WLpHAb0+NG5n+nlJXGJ7HIDWd8akVW
SYmaSbv4Yd8qMDkg5ReLsbI9JmcQ9TfsOIP08lEsqTE3S4udrzPqkH6MXRy/McCLOsYPkYdnGd6f
snh2T86pExZWL9ejIhlnCYp/Vd5umnWOxnhzT6dRSvI+giU4DA+tEqOwtp3fuk5Zod7or9F5tu1X
90AHOiR/pa0MY6WT3/qxYbnbYcB/fl9vVjY0L3gKM89p6IXFmxJ97lXg6A51rCSW3yR92SB1TjH+
lt8sI67lAaiSro22uDS9drDmHEYJJTs5uda23kU2U/HGn0CK0+1rlTRiavQvxkOHxwxJ5Zt9T/UG
qsOjKFuSp3CWtGbh4slgWGMt5f3Vi7d3R7Jn2luCxIh4UfuRCEZejnqvTqTFu5E3PSK3xDRw1Z+z
NfUevNKfnQaQu4oud5Rwx/c4Jr2u9gyxsU9OW1DeRU6uh1uh3SvC3mm8TMaHaxXvtGkvYZdURrZP
UuUUOtprWPnA7FF33epyLvnZZi75SAwMqWsTfKfO7GZpMABiZ9ZyjOxFkTXWYSFgNNL3w7ywG1CT
SBIBmfdd0DxqOAaaRVljp6lCKaE3ePlOmk3m+LIXNjWloPXnir1U40rl2x+U/67n6g9NPYc4ZJD0
4zaZS94++zqHDacSDomDgF8yaDIM4pjJx+lLuSJSFoQV//Pt2Kq3uSB+c2zy924YMy3+jroyyznQ
kuL0ZROWL0nxUkb317FqPyRlyqonWMpVm+8aHc+5Oa6nGRYzgFrNkQNaZPFOwwzDnn7kOxeD1alL
oKzYPIaWeuHpgdEiHqI2cVSm8X0tRDRX/VkNvnZjOKwwQnpka4s1mI0MPYci0/FKyOuvnu9rCXrz
uRQu5rSDuPqFpRhKWnWTy0EN5OWlMrEbzvePN3naqPVD/CFDMKR+HWO49GJ0mLLP9FZJre/uRoQ6
In41zu7rwI82mSoe6ToGHRM65mOG3Sj81TqvTvnI2TlrKrMinUtUx+eNkZ7jkvHRzOIYQJn74Fnt
mXWEYG2UHStzMwFyON8/9GNy/hYi2kob3pNmJa+d1wiNPzQsfv0A+eEQMExMjeB4nkopKBC+qMfI
zLhTcn3qQmu6I/8DSfOwZycvXy/AHJXWid7xqIsqk1tmaBvb9P6QGbZdqVvS+wTfQlgGaRLeu41n
SyAnygdIE/sE3lE82AECvmCsMYTDFTmy92nG72OQcLFC45yQcrXF80S0PagSs71B/ZAAGMoNq3LR
vDnbgp0nKPv5Ihk8t6G0qF8xyIw0DKQo+HVZm9LIIucM5KhPntolQXsXu++zE1H2Q6JaAc7n/MYe
m6EwPo4cwQzFvj+n7U98e5cA80Wl93TU1hLq3jCiy5+4g6uL0q7msEwFDSfevond9iq+QZuVgSjz
V9F8nDkHxhb6RPdoqQnVlg8tioLaRLz4kL82kDbmFP0BgwIuE/d4UNYdAXlybosxb6EQ+GZ0UR9C
5E7BXCgIdYTNT3mQA2fR1MhmQQn3OGRl6VKhRS74ebzyTa4zSTQbkyXMSVO6DbUk7XfLyAF5LmVR
yP7P0oHSRSnaxr/o96rx5wynpdSxk4dO+pSbhLGa6hOFV1EuxFwa5Ffy1mEeC5LAyDn89LHRHi1e
YOR2oZdJzH9c/RQb7/xUSvuA/5d5TbO6KlBUKgdIK579ioNm+Djo/SD3Rz/6HR8f22HpFHf+iWrN
g8mOciy635nBMaxsiHgQwBkEXkGaXhGjj3hNJnsRtMqzWrljhA+0uQpwV5HhUau22n5bdqeZ6she
YXki3/7TjvZFR0AEu4k7HNnmxyZ5mfIDy7bichAPnAYP94o/0dsGtiuPZicJFJui5uhOxnf9giij
rKtIGgjuZ7Q07PldfZE0mfJ9e9zDWKiNg0g36TDEkJFl3TACATelHwLjQ9JVTlIrvSXR7jonU2sf
rX2IAjBi87/cYm+OgbCCOcP2PITUY7yPhCyCOAZH3MigqWLh2tH/v9FgSXRsxGP3utXPlFL80eaa
Mocg5YP4JfsFwfcHwTOeCKUT4zEb+Sh2hM3bNKr5898IEKvjhJ2pPhd/3z2Y7PIvH5Qh9hZIPNLx
6XBstVhR3zg6J5hum6wEVayX4QyIIfnwROD2fFjc+p2PRtMUZQxVfu8hYeKiaI4bQG2rw0B+a+Jx
js+Q/Uekg08rL6k8Htgh2xU98qVlZ4l8ERhG00tWFk7RMqhi1K7vlhrKjhJNvI8n/dy+oxTm+RPc
u5Iyryu7HXaPDDSmGV5LiJ6OeoUsPk8wvzkDJG0gkPUAdADt5DH8NPft1Wlu8ZoWmRS9CY2nn3xK
GwmGhQGc+rrfPFkDrHDZeovKlzJqI/N4/cfTZOX3w+CNwfp+a3VnQ0SJMZaS1fKia7TD+aQ3zadb
iJLA5Fr1zWBBRhX7HR/Vjcgl/i4K1dqrptcu/9jE+2LjKS+qOY59E/DaUjZalmdg4BLBGVWar1Xz
3kJto2aXhmcUneEaImiEUorSGpAunl5Hq4SI60W/bszBUKAA6WQcH/BkkuPe9nvA08WrJAQKznTc
iHIhdTyATJG2A8wQyLSFNhNV4981sfhkLV7Nt+CdDSqVLbgWASSwPgLhrY8FmGtYQRtetMX/RJUb
tYrVFaaJaT+qoZo6vtIlRKKShojE0CJzeCMdP51Xvh5rsdZXothi/T3ybsn0bWBCs+g2KJkncs57
pNfRNSWrn8OoGD/L3nfNQ48J0MWTatJwghVHiryYOA5znt36r8xeP34Xuad2EOCt4E3pgWH9NbXA
3/QQb04Ey+faUNZVqezJKQUx5Sck6oQAdTalmWL9ox4K3E7N2cQkxKumj6y0L6RqevAp4INJC1x/
z2cdw85QDGLk7xOGo1B72xobuKVsqoTOwz7VGBipTbDujlDYjIBWYdTx2PYnzgnAYdFYVrnK9Zjz
gZO+3vWAmaImCF0+ppyHn1aC0wCh5G2yIzJSVkqq5WDeR7fSLYsovG1tPT9saNJng5axyqm4GIJT
Krt3RSKgi/P05AINZstntRg/U39Bwvtnt7OiaWavGeSwM7r1cfdRVOm3UtxGa+OnHswDDXEFhAKO
elCD70PQ/ENBzDyonR5Izm1rwvg8I1bCg5BqNH33fnOsGCKL3qjg0sA9xzDiwOrdc3RbV3k+TUhf
6a5LhJiQ+NsRLZgO2wSaXwqti8DeD02nO21Mn7iFwj9QxsLsSHr803a8TLO9tKncC/ROORXAiLTg
2yGMd34Gb67OydZKUN5wrJdfMcCgNEB9m9ksT1bBeN7As5vLvM2rNfCHbs24fkoPUiwZM8mR5Czw
4GNxVfbmj+gySTq9DfBUhz2gDnoIXF7OQrXKLz39gGh4/ohXUoAa72yaGUM/1TsU+WgWHX0D/4ro
h07zc159P4KnLw35XDXizHT4OpAMC9tmCMRVMv5cHmkoQczZRZMq0quTk0VaSks63Ab/MceiR6Ji
9+VsSFMnzYg5+KKeEmdQLzEZJjHkD0m/Fl3BYMYwJwlSp8Dzdl2+Q7Trx4R/yBZ9BMHKEWbSvWsc
qdQUYnby2JF/T1qxGSz0IQ6Ybilc62PYBlZUarznuR5QT0OLnpcO7TS0fSR8Wk4E0xhcaeWtjVN9
+G6WG1EKm0l1BNA0xOWrAWCTcOodh09C6Oun+iF2Lc26nkPJGNOVxW4c9Ug0YLagvCDfdLwd40mm
sANgNqxRzu+J2+6UeO6oWW1B/KRTuWA12a942znCznv6zu+WPqwQfX8Lgt5JBRsJ/iqh6l3JYClD
sxyFcGuTLPjNm9rZ9B6stWftUBm+c5Zel/8u82W7KJMi22hrACh9c3Ifw5vngC5NL29CWGVbWuSq
AtT/S9npBUse/cyEpch7qdImhl6fNCbWa1Jn1X9pRuieIpwl43sFRaRD8rFu/M7F+P4XDba079Ry
UbOsl4zkat9WYLJtpk81z0OkbwUeNORIrIyIHuryEmfa7TAQRTDVaduVg9mhAOWJL797uth0xKlZ
CfERTt6pMMHaSPDwVGef+z4WmupUWYaRi1QcEi9QchkcjO3xtHe5TgtAaRf2tnjEUsIoE4m4cEBO
/V2Jbp6euudYFMS+pvrJ5+B5r3jAdZDk9be78mHQy0LD5mTM/egf+f9iqpZonCUF2DQj21RPkiAc
0M9O1/1yXsFLMVnTJIH9Cp6sx/+Dt6fc9v2M5W+mQKCX7sokcu2IpwQtFR5yx43ECuRYDmPHkjqn
T0AOED8Bo/Ei1BBJQE8UQeNo9mG5gVNBlTkBa8o8i4O1LbhefRMdG3pRijn58VPNQctcF4+xmQcs
/gRLQG57kVdFeoC4hiBsV1wUSNpySFLOC7OFrtqsMPPUvZo5KIcCsx2QUihwQgIOjhBXFe6WEphp
6CKbqV68/e5FVIo6I/fCeVynyxAJzIYR1gyPJ+U4by+PmSeze1fM57tOqplRPehQREYqufdlYWYS
he7zDWIsYbwv3iSJ58ATVh2DBkqy7L/FAvS28ieVA2LEDDC8m08pTPlwYtn8dV8qK+SNIbuK6tcR
YxK+sak6GMUEY3rEKbsOB+K10VqhnpIaT373xm/PlVq/qaKxAq7659DWh30U35Rb9DmNRUWEaWe1
Euu2FE1AL7DPKjBA6u+ueF2G1UOTOBMRRnwE12vVzuKwjIijHEiDOpf9VGgNLnjIiLBFIuSAavG5
PCbuyr+RaBYh99O3ffo2O3j1i9n3PaihJG7YWXhpKO7rJuHCtoPKAuU7+WFXRiK5aiE+c7VyhSAA
54UYphKIP9GhDEX5VJWSB+GbPl5qIULytzPaf+H8aniyEpp1wXo4nFWNAdNPoB+eAMFup1/cWgP4
OAYWWkLAE0zTPwpAPa/jndQehbIiWabw3G9t/gcCymQc0HZ5edJbNhzeRARegXjMSrV9EOMFF6I0
vdC1bkcjpGJ1DYrDgAIP1zJBg+R+uqPeUvmNep7SuT9MJcYJuYSCWXHvC9fax5R6Zawg62tnGwzm
+ysePLSxVO/TEASOO1vO4dSC9MttgOUTIPBKlVzkKBbwdTcCKatC1hdQkV4D5tNFcsQ0aIZ7tOVm
/C5EwpBC0qZKWci52h5GCZ6u/uym7l8BL+ypMyWlk0kZGk01SsCOt/7n9k/1FMCh3VxQbjoXaJw+
iMsfQ6hdYMGEQbAiWgi9MFyRt2yhuRZ8ZLukNCgP47/b4jRQaF0me+9Q+7lHYZF9Jw2AvH3LjWyK
yxy3dNWJyshk0mNHAIkGlzL44aY3s0DCd3ZW1cQkUEt5ZwE3l3QUM7tNN44vJsovDAKxRnNCWsIS
uglGLmLLx2zvk1Mx7hcnEEyVdavqH0rill9fz/hdViyZf8/TaAAm4T2UwV4onpkriNLLtWdCbsFX
YHDYztE1bNV8CGUsaZcsxpdGtwCY1KmnrUYYMMRqlm1Gt/gLe5P3prT0m5r186IuRdgW/r9b4CPW
476lGaTZ93Cr0nYqT5ylhMk8A92TXqC9Q1+TwI5WnD3Bj36JGPYx6m71fwWMGTNJm9+Ra32j7ESE
rkvlHznufwtvzt8Fx9jgtm1UFCo/7dBUtWaThOraA9sQlVbVRj6cJW5Ww1exVROIaZ4OGDVVL+jk
2iRieBACwec7G661QmYw9deRSNDZlh8fjOz2ycsuEZ1eJTpbPF4oQxOXPCBko0VmMN+5PkB0vRND
Czw2q4aCmTYZcYmL/3ReFYkfR7U267SDxVjLSxZxXIfaxSNO/3R6+Iicsgl1D2K/1a02s/5KUagz
LoEqT+6B+RJtMxjRVl0nDKXZb2qYpK3VuTp0rCTiE9e5phvClnVBEhVxW2hHWYk3PLSs3PlTFwRF
xUkykxzDudj/jEdF67f7YqJc7YIZOM1deO1RJOZ+0/lLsd/M33jmQGLVZ8RKeFJXZG6qd9uqM7nd
PHpNEJPjrZj7ZXOZCQ6jYXadVfYx9JSyGurN76XFHod14q099z4vahtZj2ITYYN0JH3WL9NJautu
/SI77oOjlM1X7l75BOx7xu7zrwx4p16sdyXcjEIk/iskvIxRwuJBgBQcks6T7Wo37Id+3d0+za96
lP0tZCvk59LeFkohXB5SKSY37FeOg+RCFyrYym7IARAIxVBBxCGeMJoo6WZTkzGqwOBq6RoFPK5g
AZ6HVzNn5jFtQBxv+jBYeD+4HOzz2vvuDFtxdJtKKd0lR3Y2KxHgu/BvT5/VgZsmPFIG4VlWKFcZ
YGugvJcWw6odxNK1eqiO1u2t1TCpDwUM3K5ujnl54UhtxQkqemSJmBCVF402HJ0pSivQCAYjz1wo
A6Znxf3oFETrjfyVaELXJf4Rl2vfjcf8piArqGIoC5TAVgX4Itwq4yKz4+6KzEaqNZi6c2hhPhAa
On7L4h69uieSzpVft3MyptpM8lFtDd5vFCvJPZzfXIJR0OF5864FBx3d2M9F2Ju5cnTIranHssMy
kZFS8zQJd3kn43InOuHOYiWcLMTjB1mttTWA4DjFX1Xc9RWPhePJnUetenmsTHh8FRoY4DfjEMF/
JrqXh5Cp+O1WgbQs4Uth2Fxx0p/tIQ0Ki4IgvD/rPnd4xdhyVynMmF+3AjIWJML6Jma5x9FVVClp
4PvO5pAdTtxTDExJY1s8lsXs4yQmeGU2z1VzA+ZWYjbcZ6ZZJHG+LFV/SuUTLC4CtsFpN1WGV7EU
+APjh922G2FNez/U8RWERMck3MK1iJMRVSmFHFyDEODRwxm9KPbSw0DdftO4zpnX5FCzgakJrUfD
lmJqRYUzlZpr9WCPOjv6o4MAGQsPF9yX7mDVq/ayuper+48HCAUyzWsrZex10Uxz8m6x7KcdTl9v
r4r69pZBJRJa7eRFfDU9tdWm3TdfOH9XhD+gxCqWcNbdwR2HqBMTqogoOExqEBUsSBFSpLTaBDgF
FeGDTCNlOLWRjzfYlUYYj7Zex/i7mYAOlwY6P8HNeC4xapSfD/6A3U+zTuMgWemA9eZA91EAeVp6
8SZwr/+iJPduq8R4uFlMgu2+c2ojzv0g6awDH0yZ3PkpND0fT/3NlUnIwtTJww8vneVhHCwHvqX4
qUwFXvALUd+xqewfJo6h3qPCqqPXaMGVNjojEfgPZrsR7VI8zapebIsCPL7Cm5OuBbzNIlgQ43Rc
prjfzjNEdM4YdFd3Du/HZRAj2iGMGi0fxRgognX+RhrSb7EWM0hkqOgTnm5AhJBQJV/x4oRokQEk
S/dWBGvZFcASSma4dreq6WhCDiGc8ZKl5cFpMog5PZuFeA/ieimIv1YoVV41kF1Ua5Qo+IuqireK
yQ89H1SLkPNnGXG2FShoFbNkEV/il0Wu4b8ytnNOwoj5b5N2ut8gbKvewI2l0bGIfrOWQZG82YA6
f9STSfPxzGJogYK2Crdjpwth+HsatoqsjmyP/ylbUThmPG+luo1auRPM2Iu1hHMNo4niw4iuCdgE
Mlhv9m3s7tPo//1j62orbD2Pp8gDpFLuTUXHe/JunR/ye4QWnr6ONDl7irh8cWXkPzKab0GOjY5a
rTvzoPc/QuN/YotFL8CjHHNwIEX+M+9tzHDynfVtxbVCKzgTrwuFBrlUNM0lpZ4UdruTxn7+PTIO
KENtF5PfRUpHBoFWlo/MyDoo+U2thcKQGfEfp12nI4QUffNQogZcFuANKa2n7VOWeJoOPAw821/D
pvejsKUFtNwA/8pndlKFRE+EMDPEBs1D5W2nmW2oNMP6tUi0t+hYSfVIqj6+qQIB8nFWWGIJR4r5
UmunSVM0Nybe7kFH9sm0Vwqh9JcLcblSdL9gkRWqPjmLXU/9RDr/yDOzIPDTJnnq/2LXA0XenOrw
MMYol3f3SDfivuB7GesLnENXnjFpGWGuvh4zJfhdZme6B5EbBXq3/MzkVD4Cdl7E4TbV4/oN+H4t
92uT7J/oUmkqL3v+265YGRIywlRpiQ5tMa5zo8sqnmjKz19+v/ZV51r1jdS6jYY5En2nKySySqvp
M1emLUrzdR29culRgKyKKQLtYptKtMPxRvMu3WMToVGs5TBs1U7q8Nb4y3ac8Wiy3kehZmCJmVCW
HAy4CmSzu6rA3UY4Tx6kPnoyHoqZltU+HFivo+XqqI3sbVSlviU4MSPOF65pketEG+5OEL0S08du
tDazkKcpz6AjV49awM7PqAAM5JLUI0F3LDj2yR9amqBJUaCqF5mKr2eFlnR6tCREaDRzZN2+LgmH
S79kMsdps+k4bVTA7tcrYJ8BqHwS63hKvO4VPRJxwnzPenR1wtGDD1bywOnSr1SNItsM89SVmAmi
+Yr6nj9a3gAqN/ugkMdUw3Rg7g3gD4R1/bDdIkbF6zUxb5V4vn5Cu0PuE9FnZcRkh0LrXWrXQtXF
qd7qUBlNiKn7U1DfPB6s2J1IdMg+F2fOxRar6CBAb6y7RJpsLX0vuCJo8+P3qPA/v688dNvI7fyw
RP10dKo+Swz3k1C8rwXqE9GjJN+jSDUhoJBrrk+jyc+9qOQfr7BPR8Qh4NPzgAj2znbEcmAfMVyh
lvMeAP0DPsL9jz2CBx83QaV8oGAjlRpmD5xTx0AfZHu+sYvX5uL9++i9rwx2VFOrNokRv2qlS3YM
O8UNG2RxAh+VmsLnsHrvS5R9QQemdxU1VuYhCUxgoe3tXWgSVuN/gl19Vj9degbzvSHsKTbfl65r
JnwbaVWd6FWRXXnpacjZ3DmDLOa0mfwYb+6PLk8wJKl0L8Z+X5QhgxmOTlPwiOcktMM4mYiRoAMH
TxR96ZlvGq9NlJP7U7+9qkj8fW6euA+tXfw/Jq1KaHZ5VPWdpb8KKGmy4Y2yMR0mNd+XrvXV1JD5
2Vs1LwgzeXwhY2JJ7mZz7W0SkwVazIGQiLw4M2gP/krCIpBhxhnDmwUu24os+PXx7RJhH0AJ4cgJ
42wbx30SoWDtHdsIVSSnAOlTKLHs0B0QV6RCmSyLYZHZVSBwgFR1OgYuwwmzFJ53sbwDfh+58TiL
p/MJ27HIlIlJulPjfAofhjVyJsXW1SjBr+JvVxC4XdVyGx42e4OkVF9lHLAiJXz8Zv5JwpQ9qMK5
ZFX3TqvQeMzVYkjS7ZuKljzaRCfORCONbacXOYa6SqQw656XjzcQKRprUjluwCXxnPwLvEahhiZo
wrB3aHuTiyonxIvonTZTrVw7xLIDtyDeaI5lkdtBScZdhaTWsskKH9M3tN6AbMbZHQMkWxwkC9xl
HYX2stq+i7WW/518Em+xNSgHlTvcdbwZ9Po8Z6xQVKNWd+9PB6Z81encrFKgd+MXTwJ37D4diReS
Dw0DLfg+G83J3QUGtrJZ2vIHYSNNGVgCyYRLju+YCsS4Bp8Q144LIH5l89WNC6NXiRJjfUq22nXj
7uiDyjc+oo4D+1llMs0aia4flGqRt137pMwsRxGhPFAq2eh73x6sN+iPT/fV+zRzcbdDBNLeTyEO
/Dnw0MSHhBJbK8oeeDn5sh4o3h1oHG6xT/EjfyBJ3D0rsN9ADMc32pLLkQp6FeORRLk+YtpvDpnA
KgfIG7Pq3ne8WEQqfMTPaOkLYOy/T/9RwcMsem2kKzPwldqgooN7YuKX6HUWChe2otSdb3gMOAMr
yw6Bnvxlzp4L/uBOYTRtfVsWikwDE/VuHBI3uZ3iQDTUJv+q093RC/Up6mMDggrfXg2mwZZdqzor
zQHcAQmyStb847KEtqgdJ3ailOr1Bq8eGtqJi0OVfvfhx2EROh+FbzYaI6RBPYlHA+eJkTzatZIg
ip6q+o/5qdUOV326j1rXXnMbC50D+VMpb7tGQP1G8ItJ/NJe6zbXT0dFM/J0EySAIgc2DN+z5aQX
TpjPW6hOpcnL/KpginDLWtYMSc5wj1psdab1Gtexp2VEGapxOmPcxy/Zkar+3QAsm/QdKNBh7Vvx
SLOhP87SiACuB+1yMBtRAcbqUsRxbaHezY6pvAVl2j2qAS+lQEQC9ZBuSf9tcbbVX3MsZPaVlVsB
OpwkdI0/bUv4U3QIFFoWf5f5zlsaz/7VOqbafI2AZj72IdpPp+eriEQ6YEc1lqP3prNY3kQr5rHn
Ppb0NBrAHReqPqnWqgly42XqzCW2YyYpHXsi1OybFL5j8Y2s5np9NflFxiOxOIAyDscOtvfBq8XK
amlV0JvNMJBieavzjeMueTmPLYQQiHZlnLfjIdc/XZsbHMkUQlr/qp/IdQsEUGz3yCPq9EY08hbi
UCdx3kRBnLB6lEQ7YMID0OBNJEe4bdOu+bD8cUCRcWkRI6CJ2wmmIN87/vPIJ07h+Ab0po9ZwGkd
QElmCnH7fj0unIeHLN3AGNXmpr8OhCJH7b4f5zzmhW4GtzB2mmUQE1V4HkfE7dYqUh+IzuRCRMj7
SkWcOO37epoRZtBG6zgMEXVecPhfAxzgd02BbwMRAnDaOt42Q2HdPcy7B2YfMiVpOmhLV9H+jkuE
rJl4tS/7M1gpth2ERneMXZ+QxswijEV8ASV0jGDYTU4kwn6zVU67ReQT+iogCf91ILrwPGqRN4AE
joG8Xjki2eihhLP6u/WN+qT3s59PJXkSOFHXWdZdjAdaPirxAGyEw6mxtTMics79LZfGmcqCbazV
SDNlt/L2BK3d9L965fxyK6awZ6ouERz7fZTsUfQm1Z/bQz5UleWakNHhs2ablmN2EbDgTk5XKdjl
bChluvT0bVtMat0nCUVODPSUhs2uZk/38XIvKdcVYEFcVkZkFjp82iM1QSuAk+x3qc1YvZYMzSkW
BT9R0ZEXni170W/f89E3b/XJLrpXiOMkp/pbyDg8LVqGR4nPqAB15k3sTBjn9nav8oCYiYFENJ55
v1JXuf7AMOlGedxjqyg44jSUbLTlkQK+rBFfdGwj6HB7bebpMUpYUgexKDuDM9/Sa5wp5SNN8qXw
c+ZEN2lwegRYvx3iSYWBErCJbVI0tcANuCvH/8odHIhLc/6wLjEcoWD1TJ9sZbq9Ln/20yBbLXi2
ZCPloBmGGg3/iES7Wd4dmi/cDsiv2WxjNSoTXAfITUUv2t+idMMmDA2pccq9TJ4HH/OPZcUerqar
XOHyjgLO3K5wALno8HoCzlz0xPzbRGyMNHMtlWNH0iU2n7KDF31AEBPRiKpAaYQ79GKz8mkDVg2f
MmaSdYXpE3aurzDMyK6nAczSJtv6A+pXMgicgl/WL19JuyrdxdI4WwIQUym92JcZZuTZoaJiAoEp
sj7OQfsyCDfIYp2YMSiF2KgC2F8y3ir52nIXw6L2a+hNP564FP8oNzHo/nRQEy7Zq17gk2pXLLU4
9y7VQNMtGhzpTQq7nIAtA6S4jm9p64iOgTebS6qCL6XUfDzx/3XXq1AutFfwct7p2AD4a9LyFWiW
Xy/eP1mMoADlz0sbZioD23uUuCOtlQIT/JIDna1SP8cQdRMuvkpJdo1TTZQDpqhk3hZL/LozOKNt
974Fe0VWAjQpSYMPbtnK0lsspWwrdnsUJ4mBD/ds7nnqG2akRdAd25guiuCjF3PdcrcImkmd4H0i
MmpSJXzAi/UfuXNdq/xt7hKjzFb4msNeE8RtFey6oBOZNjVSFt+gfP0qNR6fmjBZ0PHiPMFBxhSo
HmDZoFVgjlBgnVnZQzdmgDFwHv8Kjct6hKMTY2pY6EvJETOsYDXBgBfJ4gquooc7JcVGdXhepgxg
0lr7jsgQBru33sqjqOSACqEBvTMhgC0fkH9FGVD6DEDsB7U1lSpmZm4zxTSFYH8m+84lGhGdHW+X
r3U7esmUmS9M0D3XfK2U9jU/ParkK7zT0nN0WlZnzlgB4V2+MxF4dq9u+FIua7dOmiRrGFCkpHMO
ChUUaa7kE+K+7SEPJQgE/iXsdhTrZfxyErkgTwkW7c9XSooWzyZxIE+pKyR4cmaHh9S+vaggXLQk
hVjXx0mQ6Pi6yl3L4ShUAZaNlzjH545YXGg+n2Wapl2xQcWdLVbswsru7Cspqe7dDkLExmQa4Si3
2xnhPlHR+medCEIb7nbFiSqPUMSQPtw7AQmEIngj8bX5CIab6V7uZYfN0/GLXN/6sR5mc//Y+Nh2
qwQcCi88iSdPmfi97z9leGmyyzSbcrjcPW/efMPIP9WqdxOLCydS+9vEP0TvcnZB78LoUXStdCUk
NZ42NS74+wwkp9YSlVjJxJKmmTC7ogQsm+uQB+pRsqrFASnQIPghf/3H06BbgQcNBLyQJB49KTj0
OBl/MTHFPLbEAmJlOFz7iL3KsC/gj1eTfy11FTp9euN0XPsBsqmXGLkMnzrcYMN0Jeg5imHRZfoy
oPH7KEB42vr5odeeI3Cq2Yt2nEVjiShmX5lBP52WItPFU4K174l9yfKfiujnudAfrqUEAzc1igI5
D2k1I0CfwL0rX0u7OuktxJEryzK06j+d1rr7oaNqO9abdMQX7hisvnthLEPSlcjfDNuPjw3ZDP5q
ZKDoudweAHvm8YyNCaokmPcI/ticqFIe/fz9aMgoj+wa6vTb5+kY80cxhysqvnRVIMyw30u3A3IB
c+8Z9n51zzm8Rwgtmw/2YynYznUmUenbMSEoxCjUJ0ojS8O1pPZ/racezK+2mNuqvxwX7NRfo1bp
k6YWIl+SangPf8KXC0q9jNBOIhloaYBsQeDvYMlBxUsbpUDOpZ0BmBpTtZ6mW+peJezJ1NPxWi3b
LpgZSpv32WCdaCMzU+ztFOCX6907nm8QopbCx0ItKZjZRZxb6wHv6vFCGD5AiBY3YlEmK/xzRBcm
sZcBsuIbFuJTcZLenz1zTSoJ/K46c5PSTAnwsykA/7IAnEmuOcaFGCaB3WKIVCEc/ax33jUIfzsb
NN23rYeAVN9vkFkKA5GBBmB9hCxjno0NInQMMZWQzxcgpo8NBw4Drs5rJtOn44Iq56NfzDYZh4Re
OMUOv7E3gWVxMOWbQzfUtCsjosd+m76aYOJb9Acw3n3A3VsPbb88w0soRZ0GE4pkQJBwJSF0V82o
KBhjWWMIqCvDiQYLu6vq5VM7RNmw6KzCxva47T0JMGb7GEdc+ccDINTXo3JbTKtjro4nFhvNZuzl
2FtXnkSmU3z46LX15prfF5WdjfPeOe4SGnGdgQkjLXzE9egGPuGqBHpw42mtsW49pbUEgH9X4i4k
jtn/SVCOLepzXFk7n08HbJV3zA8m27zovOXoNoa389Ovxlo+q5pwYSFK6VAvR66JPsnX114/1ijO
xUOPzVIhThRU30r+pobHiYw/0Y+7fI+afXrX7cHTsYxWxHFnnuXAkqVTpJzMHLDVYxK+sxYzC1jO
tVH3yG8tZE1o3wF6UdxadaI/H2oorpaTS+X/ewVBGj8xPlBEQUkfkkgNKhipU6uT4JbFuyOrsJE6
t1xJLFZ3HkNbN6m1YpVanMJBlO44uTQso4Q2diDDkc40hPZrHlbYgn9W6PVgvWZrpjBdhsCQemvL
X230QnBIiotVsJqQHN/5Cae7u7PQTP0GFJNvFacorwDttUvVPwPzbNUcCkDIlLSN+AVToXCorjY4
uZ1t8pbrWGJVVJss/o3O+CL6dsxrb+sARJjYgeNxmY82XfQPrSYUpsUz2PIH6TxMNelmjMgMN04p
iFMW/hWhUO7rQhSecki96F78flNMJ3ahSxusTRigRJpPzeRzGuyWi1bL8srbckkl9zcEM2SsDe7M
6vIZfIOTDfedpu11xr/nk5dNypfOh2pkIinxaG8o67ml02OdOLknmeymZMnGOIGjP72ECkpfwHB+
/SUsor3fEFFWxSZZnU+gphXi1D0WCHZyFaBUFjQlswyPGT2T5fgj7a+7gJmx3eO1Xqx7huhyIaLT
E1D5GriGuDcjtngQbJSVoTOOTh4BU+013qVCduGJF8T5uYrv8rA5qDO16+QfSCdrmIe1cYMfKd5d
62XxCpquEJq9rSj9XwxNRNC6NpqBm+R41cAfqaPawE5uRokleGny17niMQWBX2xo+TEiEFqApusW
jhzZQ5X/kohQWsd+0kVJ+Uc9gPGkzcBV8uecYNOxgA4Ca7n9dbqbRYC2D5wZ4IPXe5cuBRqmRqv2
1l2tSxfkmsDFgyiqqV4lAOivBWdARRVmL8ZrLFjYfdzgL42Lqgl1/5jXI2l/+PkAao5c4dWBV/+b
cLltZy3sUnAgLM1fx4K7CdwHsqtyhaJjTqetsDQAWbuTzAuM3AmtwWmhMjdpgxfkSK6g3EJXoTIM
flul1ZgcFokuaoOvo0c/bIKDo+4RMtArTWaR4qsIzHfWuH+X/VyrgtYrinwpYMjPmNbFTAhNBQ7j
qe6D23ENF92e35JUBWxdSvfkb38FQ9gp2JUCxGrxrtqaJZJjKC8QBj+QV+luwuOmlgjFe9Iy/xf2
Vv/jFQB7DQf//2jLrB8rLrZZfe/mg3CPj8UEAyyUDAyi2/VsCfrm35z8VCi2V4zY9ElfWzdBN/10
fW8KNrRsUr1bjaPMGTPNIjZVbcBFArAu2N1eLbWxIGG/IyooOe1bjslnugK6b4Y5dpedET/jEaeu
kf5+bu4lAoKtuKfi3sdyj2OYMCpYolhzTnkPoHcdQ+9VBIIHcfmBwRX4+4rH4C9Pq1fu8D9rp3Pf
W021UhvIYd2TZTfRyZVkyDa663sFMHoQuln02Pfc6I8l2IJMu+GB8z3/gsIxboLDEhejrSyPfApG
aS+cAWN3F6Wm9019DDb2kqEpO8lKGpBNECd/nsQ3+5qyNueDVmtPpgMA3N/QI8C8BHE38IzD53Y6
FrijG6H6EhzXOzjhdcZxjhVe7zxsnRZuk0tOPWNwA6IKC2Fpa/ogsgqh2l1Y3YiNWaR3s7k56YBE
uM89JdaFJ3enmySEldjf7FiqTYb5i6QKfTRN6e5As2d7WPDIDX3tdeKWt0t4t82ltlfUmwDuLr5e
mqpfxkWs06+81T2OchpwywJmCvXa2AQhExSx+HLwr/lQUjTDHOBmXRgUYaNoKaIQqycsrPom0WEe
ZE+jKDJfHTJkK3mATFfRNZIeFEILFjDJIaIC6g2fbvI9X2V2S99+Ad9RK15ug/ulIm1EGWmw9uM6
CrsDuM0nzAXOdexlFXlyXFQRSyZp+1YR24HEweigoUdv6vw/ssqlL7nVenKnKO1ohNXIdAHjvf3c
PPvOKraq+sTFOWv/aJsEJOzglX6cLjB9sY5dVA/k+e2avmUHO6G9Rpn1KGNma3qEep6VNz1o6QLB
ZUUBwKfeC+SwTQm37+70ycgGyGC+DIsYggBZfyZy/25w5HJPeG2q/i1PgA9XffbwO3PR0Cxt8JqK
P4jk4z70B5u3q9/U3yyHQrdNpxsb84vkFIyVVZmJzyt6t4bMm6KhxNUmeRYV+hhmqCZHSAwTssGq
F74QrA2T97XTqCI+OkVXBqKtCSe1opHTMZtd414pxfEiIuYHEO08UilBGJD1N3KLLJnzUbxUwRD9
EtTcx+vdjw+oPx1oRAIxqXPw6byB72lJdbeuIBPV3feZVOOdVTlVgB3qvqUkWruqbIIevIXQFAc5
umQ8rhOolmrUjU60Ia733ccXkl6sVVdNmjOvSZW0Dj3VZKSQe80l1dm37vBAOF6HwRsGw089oJ0P
d5wNu+oIYJv6b/bqTo/C4HhYnQhk+b4wUeaYUAVrlnzSu7INCPVJS+9FUi1FPukbEuupC9n/kLoi
IyFVx5s9NiDPdlUwOvQT+FLjImD/3WuD0kYdUTlTrIvxkGSADVbns62PL3nHsmDZVX+7sHQ5eA+N
6E6P69odOzBIe3x7nG7MmHXr5PEIxfX4lF/BqnEJ9hy+TM+oiSjGi3p23liF2aEwBT+GxrjtVRXW
6O2lNp8h5ClCd47HUeyQlyL9MDSgF6b0JYWux29FgWpAPBxuEkijSTfAR6p+33eMekUCS2RA9IFO
BEOt3n//zyJc3L+W94Tgo3nRR62vRTKlxQuwBe1CY+u/oau+PoQBqYvkupB+fv7kEIsFXR6qlAUz
UtPbsqVp4gSE46kdQqm5UuOcSAG7EdTpYNSJM2rP0yzyC5cMMQTPW7hujxX1vY1Yr6TIhBNa+zOd
/8m7xIQN81VwtdMYIAhtbacgeUODrsZKn4PJbiIj8bNa3VHzvC0sj9UfVN/zi0HFVR4QEgoKEAYu
wB0vu3Ud+OvpFgiojaheRzGDmmDJ4u0riazR8RPK1B+ucJ9XRsNqXhMc9RusL1TE5peNxU73iESS
T+BNGrytNQ/8nFlmXlYqZ57qz8no2fIQmaAvc2Vr18H63Epurmrn8LlF/hryjOkO7cHpmqIft5ZR
S0dWBgGsPJrIwMNE+slzAR0JUf9WDFAqUELeEiCPXv1k0sYQ2wF3CBpWROKeUSmpLWx5KmNOFOTB
cpcugIZo0jf3km+Dati0pti7CQurR56U7DVsXs4u2xoOQxpj991Lsxpi72Guwl23eJyQh4tz0ANC
ZGoJCkFNbSyKRYjB2c48EF10VAgfxv6kGwmnP7SdJATJS9E4FVk879q5HeD6xUcloQ373uRzFc5U
+kAIk0aXC/Hokp4rbZBhKCujiZ/za9W6IKyb3hVs3cTeOT33ED4SUulsyrvbvaQPgoCRIs9orV+z
t8BinpVkGGZAXsQgpJCA3TCX6D/xD60xIfaaKeFuhRJPUJOu0QUrBfcIuzdIubw+o4sktxe1dnZu
4vtOkOODKjkHhfNrjO+mT/OYuDgg6TcfZcovGoKw9UO5fxuAPX0jSSygeaO5UPqpH/sIce0qyJrR
R+ihF0coH1y3cDWI5BlXwk1yXgJSDONZQOwV+2nq7t2991OBymUyRLDzx71oqbLu66tNd40uKL31
OwLX+vCmky9b4uIIaWM+7qrF0XtrAUI1ZmhHcc/Nu+pqgAfhKa617yBCVZlfChf9vxny3MXAelHV
YYEIy5Llh47Y9NExvITI7GUuWPLPJxk+VqvsY6/EiiPwgnUz7iMOAx8SHKNoVV1pZdshYiak49sR
6qE4K2kFEHmHwdCKZIWO0iUO02gI7LIa6lI+Qf8corGUBfUfng/tD3ATFxkHHuJKWrKsJChESUZa
A6JRzgPLaqStk26deQaja6oNOw3s0fHdDm7G7qPZ9bj5OMFfrehRrzJv+CtkPReohIVp4PZ6a+Mw
KePTI0BF2hEyHAGdqznXHHrvt9+GPD9CLyqzyOmFUGX4K1lssBAfZ8U1NEbfcoezQVZ12BOu9Y0g
Wmjc2femsRBFx+ZwOKKXrVrkLQDgKF1CovafPl1VTHvECJbnDvg20FZGeMsHa/HT/lKcgGePXodg
zdygSwleeRhbW6VraphsvIPvSvvv2v5Bv+P80+TgGdAqxbO0QdAALfmy7hiny2pJUdj6XUndYUO2
lbwVUC2A/sV1SBxLgiHnrQdKlY9jRHKxHfCsItEjj7etTJnKcO0HmFTe098TH/FqxxheRomYNrvO
atWiWcMfV70cqfJpi73WYjRCSTWgP7lNehNQRHvC8gDITquAGwDdpUoWA7c1FUzZ70VF5LjS1Zx6
wJkvAC2JrMgf6QAmZNEsIVpvJxSNu7xmUWbAPp9KMEpd2FvIWQ+VDObPhNiTCN2h26xnjY1btNom
zADuXJHsn60I79h8kTouTpQ++gUQcYQNRsKd5d60PrRqs47K4Kfjk3vN4pO6r+yA9WPML1SqyIdL
ZY3YvkePNY6IpJ8SFI2sDYle81elVB1LVd3LYln3I9qzF8mmQyFhVwi3ud7uISt1J+MZEJiHqoFM
nmnX2Oop+E2QnMLm8XjkKABSgQHkn/+60oi0Q5i9yeEqT35+GnUNIr0G2jMj/xScdbIIzrVdvIac
W1xXd5zVu3wkD6MbUX1Chak1amd2MJI4cWsagWMg3ij2Wezq8yLrejzKj1ucQSdDPDSSISvOWr3w
ymfGHuRXSs4VVVD9txCvfjiwAs8Q310o7jllv/Dty9ujmd2Vw/jNtp6mcU0l3hkcUyH4WA7u8wFP
VXGWHt/iq8fXevARJnns7MVzu12Mt4LXT+GHTWQSbTNekv/8oBCFAPj1EdB37Q3RMSzYm2nS/QKN
VcmK6+XdwD1ncRs0XVT2v83lSVZwIn3vCu23YiaeXcCtfnkxYqtLpT4IDsqJNsK4gwltRZcKgNCK
BJDrVqyiI2+dNo0AvjATlMV24gqIGYs8xjy+V9JiT37e1CEsvGBXFZIaulJH74I6gamsT1dG2WPA
C8mwmZiLwu5nPSqJGteFdNgs9pNSQ8tLagEynJXRJxRJR4zxIj3yH9m5TQbSfereoXENr3IJD9Uh
JzTskWiHQhKJuotNzb+bkAlNZWzwlmOJMAvqp6X7tbka0RtTDd2WzangYRKnSIxtb2lJ7NsZJiA9
GGMM0BHU/ndmTbYkedJxC/RwIWtIv2OKP8dgCT1QhZpqxSk00ciDs0uTJbnCpK0c2REgFr6FEHKm
mPeRcbBd5YOS4/O4H52dMFlKQrvFT/Ns5nLxOaeU3cFQVLbCO7oLEeM/VlZe0wDubbcyCe2+TB+c
ay6zwE8Y/HEURqpZiwYmn5fkZIGW21Uoe3O9asudWLBmdKVlWnzev5rnjRZaiGQRPrs/nfma5mzP
XaYbD9QXJTiPB2q/jbQM3/2taOGJ2+uAgrk0I073deZEjvPOwl7lQ4Z0U4RIYwH5P6t4nuNrbWpD
539ZZRRpecCVq7rPcFgNld2MO+u+ROeFOdmmBiRdON4D3+JbO0i+OXTjpkVQCZvYhXHGr8tXVdFj
8gzTQQ71cvTvlbxorHtpKsklmu8Ntzu1MIrxD15b2n5jMf2MpmTDEYJVhJSOYOZJZL+nnbkdIJXq
erUsl/eXdycQW2MvffwL8Ci5F0QnTL3mua/NET78hHsvPMRTbMG1YMJu3IBr6p8S+NcVlQKNjRtk
nvsDETG7M8x8aebks1joYEkMVT+TeI777nXaq50qnaFuVPRdVJw+lJ5GU5G6fF9mGnpM5vd+ytAL
kPke6NYNdKtvSXvYy4QUbmEpmjmwFR8xro6gv92x3HbWY0bH7Piv0hkHmJqlGIp9H4/logwDBLsN
eyU/2V2KfxAyfjvWceANJubBqRi5NKneqfscr7GOzZadrhAOT47CZUOaXjAzuYWv5SiIcw8cwD49
sj3x4Sa2Lh+rUllcSEBbthbr0yHveXCUaMXQHF5RJk2CIQ2dRP1f5CAxqrxvAf5a5PVwx3qbur2e
UR448qeWxv1x2fEyctzu6E5yJ5swUINmGXspJjBLe0QFXYj6P0MqaWyGuZ5mo3zGBwWPyNlVNT1G
+swGDXGf8MFWof5vhtzxZNZh0/ETsA9Xp43w0LPKPiUFZarxxYDloan6igDiRACMKSSKd05CQl8O
3rq/1hBW395cB+NomwiVMhd7CjM0oVnUZ7TqHGUtkIFDh/iRm8VoeJIYcbjlSfA28PS7kEe/sII8
jinwXkXs3FjQK2RYUs+wC5hm4ri9XrgvqfjvuGG220UXIYra2ZehiS+vGD9Pq5KclcN4GAkXal3Q
eMt+ZD3HL9YkQ6QFr7/hnnhUbjoD1oy55upU6gPrxF6qpZZ3xH+8t6NPa65o3F+veQJm4Nzw/hrn
3ZSzc8f5PQDgr9EwsEUnJacsdsCCk5uGl9mv62uLuL3R8bhUYz1ZR2prmtCkPJs9+l0eJXax5rk+
puiGEY5G8+xw3uCphmdeKufupTHLnDKcIri81F0MghWZiA8kn+YYlRsTk3cRECJf0H7VpvVECk44
rUSV+2yEQhRMEToiD/zC75tIRPjs4jkKKrbV9vmZNGYeAGmtWdQBBqynuadqXcXmbXXd/t2EMgQZ
zfbjVlZ24InyZh0aGBvZAUPFJFY45RdIqIPiIT1bRTMHW+psoWSIFh+jtiPl3XP3IX7usPo7XJLc
gHijhwzwvtEr17c9fxyDV4z2BohEgWrRwbWLEe7vLP6VsXbJr8jPkAmyPZmjGbi1SSj6iic5TZc2
aB6pl62iiIE7DKu/RVT59hrTSYexuDblFLDPCQdy7LEMBRLHw84a9WZ5Y15Spb/BBNm7E13Tp37t
grZig9QO8LUf7Bj5aMpjqSz4gloD0h0AXRDBVJiQFewAQYGCc+mQsUu6pClCJDKMAONePV9cppyR
66RfOX4pFFLpoUmioIEupzE8Juv2q6MBsmJw9m9gIhrVLA9Jvv7jKKR6jpTtaJzoKmuA00w9KWhn
nKagHxiy7IjgaOHa65qHwhh4cQMINISnmU895h89ioyrbqznBNhJFf0f3xGGCL/ymBCplDaOYY8S
ymEIWCevJuRgJHuANG8jTdpB5ERMSPM3rdOD+mqweNrotqBcWT1KrF3EnWXNLPi8Mx7tsFVOv/gU
3ohz4eyXDcRIu9/rXcs94oPkSWUnYsM0oPV8Z5AH6UBXswt5FDtgobRvEmDAsKjWFZnz0l/zWcuj
3ynvmmdbhhqFcWABbSpfP5vg3P3kprSlL0cFTYM0LVLDgQcv+DbPmEMzClNrD3VumGfbckKYCXJq
Kr4fUsn/AuM5lMFM8rr5SpzEyUx3lOMKLylDs4HpA6W/wixTla3JRfnSykNmYCceP815a+rIPjxc
1cHiFd+nDxkCYZnyqi+Ql/jw6UWvfXpTYoVHrvZPtD7RJ92hxcnfIfe8cdAlGZmsr/23lBvpvGgl
VLCj+enFzoqVwjsdkIr2zCFqZliOv3jyp7bzpQZVFlF4COKLmAeyJtCDEChFaIk/1fvbvjerJOxs
jBs06L1Z+E6L9nxqBBFnGtoppCQtGZKyBkuZBiY7bf3+ahoC5UvDOZNAuyzX/qD3x9MpggDb9alP
LV/Wy4xycQt6/viTA0bYm+y9HLu5QMIKuct2QRdzUAzG2Xcop0/HIEZ6It6K1RRXXXDyjF8UUjsM
cdn9YiZw96sRzGued74/rsswr2tofauZI0zgq4+Vw3BNPOvUPEwleArFjKN0j7pOOBK1MzmI0qT8
JE1aINKQ+hBRMoAVt7GWf5kvdlaGk5ZZ0+9JN+BbRR9HDSzD/cUaDdE2X1HkedbKQA3D65vTm54p
1Ocsm2dadluCVrKm8A6t7//XCdp/QOQmtvHBFUrYo7Iiot1FhKJwcQgz6DnFXvhKQs5V9wExJp3G
QWtYw0Qgbe6WaKjsVK8jqXSKTKadM8Yhx0Oc0Zoec8B/gUMfxLTuameG3/E0Wn/gOMNUXHP3T/jU
E3Qlz5ZziNRlccjp6SwPPBcV8RhJx0ETnU+LQXn3Ny9R/jas5qMTds0r35hhkfEFbO6RBvuujvUM
I0kpnZFVYSKAdKtNgBj0Mk9KS6zc3UXq2OiLVfPA13b41qCQGi9+tgUrI1kmIHziS9lnBYfCYFWz
ZBnqk60rBNqS4Gpn34M2g+0mLfUdZBQjNXN1dYk+RVjVkxQKzHtLtfUnRyPdkBrmb6PPCbHgEedr
LgV58fNKaOhxlS+kzfbWnnVXVNjSlWwpYJYbifITpLJF9iOLnQz1U+hAMCdlbgG2AHjd8slUJlTx
Dvn5tE/CzAf/a3RWQ4TFwPRSX03jNlqJupiUDpNPGTkcefbCFaMm35oymW3N8acmxpKvy++pROw/
p6k6ByVD+lxkyum1LdWDSeXDOMbc/pMjtSgVFCNX3VeSH2t1MfaHBylG70C4pK33RlY3aBQHTPbH
K7MZ2WYwBmV/V3Z9kEYHh+PLK975s6ceyD0hUGrpp5/ohrt5JLcwMQpdXgEtOfblj1a2PWQbs8lX
RfyYg1+GvM/Ued4A71ZFsNC5LZfKqsq9ply2szZefajfoDsiz9IfraVTcpI1fK8D0P6GwXmtGRub
WG+XbgZfOZEkvTQy7eJxLGpPgeiLFr5NhzPnxODr04H+GYEcYu9mEIZFLjPWVXZiJ4aiftavmGbA
OZZ0wUz/ZDRM3T4OTYhVSwAcOl5hV1/VIsNMirSqc0XufTJ42es2kYzSZaYMAF0jtyeQcm/SxtgW
SRW1pEJ4fKMp3220Q20oWSWrUatcT0PnKm1sHAufIO8JQ8nbXyPsMZwq3jHhu4joRMaXeK3mn1r9
w62dpibV6L9eSCN426FMOe7zIAH6b91RjxQJysNwWKPFih5BK3kS37bkBJ9GS/EEw/ryWFRQJkp0
wT7IBO870FT7vjI8XhJrhGlfBaGaZnlOgC88H1VH2zIfhPYHPorJ2lg82ls4xzzZdFa8hQvdeVwt
jh1+sAqz+6DI0pf563+PFZYe1W2+Q4+bAIoPtwgt9Ntm10K3FP+l/a8BTOVu2Atmo0ZELRDazm1U
tj7RcPBjeS4vaFzov3gSfXI2uLOOf9dlKryP/kPa3zHfT/JVWx3nBfFY0/SSKJdLj5qi1ZI6iUZo
mBSfYoFG/fu+7w5y+gys0a59FzUpYZ6TedxxufEWFBM/6hCflLvjkf4+zWZMgetwKlTt85ZMBoym
Ixchij783f7YCNmEwpCpodlJg/zaEc6iO5QzL7raHPcoU3E+EYDJukv/cRJ1SeeM0QkeXHwkbpoa
/dIo9CBYEq2rLOw8TP+DMNOUSf0V0T+6WMVZAG992hsu8uuwQ4OCn0kZKvxuvsXhQ+6bKxWGwmiz
QUwFBn/5T9njXDU/HtcskxWLUQ9wKJthUDm6JTAPhVj2l/uU1NXaJIpI/6IskP6O3XqNCAuq4p6s
hSBijNagCWTCvyoctKAAjhGaC5+8VMG7fatYNvfj7FlaRZkGNnSGk4tOAPX0KEs/J1FstpBmtqsJ
VJMmUdIWDs1uKHhUFMpZ5mMmQkIqJxvzY6/KL3m5hBLDKg8SgeV+uzD+NvZ1/nX+2w/toKJbOzUt
9Mg9nvtNeohEzVjKCeikSUTjxyiey27LN9NoBhjiw9WTePYUaS7JHmDxp2uCyMNFGz5DwRZZ8rgA
5E/IOJI91XXpzcQYvxkugCh8m0dn6RDqZxmCTWyOcLmWT+TcThydcj5oX1wjAPst0Y5PFWqwvNfx
Fvwtsl9D5bztnxjUeawsq9aYrAD7o0sIQlBHwXj/1V8A/iqjj3l6+8trrHPuywNk/9AZUvShgGFF
NOk2nnAagiR5ceBUUCuUPV9RH7WIUlCeRkringmWEI139qT4mTsHNSHk+yC9yCO6vMSReLB36YBw
8i6ZLWN5zhVreFJXAZdv4VoVdXI4JH1hZ1l4m9BnIXytZ0NlW2RStnrS1oyZB9tixrWXWc7qpOCd
UZMNfkl3O2Yf5PJN4/ZjUTXCBAUdbjORJXcilg8jjA/7e8H/nk3sdKLeOUekQuwtxnjNNpJxESvN
Qh5wDd4rFzmdhjng5whUATzCFBVtct/0rGBnsL1Hur1NQRczh6OUMiQzaa1/X3JBL81N1iNqMD+j
9D6EM6eqJ9ooDndN2xZwCCeaKMTcqLfAnQnCqLaie4gqdM/3yRF3XODkOrQ5L7rS9oEk7M50A9+M
13Clmw2ef3U5Gn4j1gzQ6Zjo2l36CDWu/bchG+cH2usjcTsQl7ZGG958h1lU6SysOidYWNjWDIKS
KH0jRpZLLUGoufsqIKxjSB30kZ/joPAyqEKYZZHVznM01WakaygSxjrDTH739c+qqUwW+wOeF50C
bgaqVrkkEop30kIH6eWTE1F+Z83IeFNWy/GOf0KLxld8qQbd6S5+Q9aohYkOucwhBFLyzfb1ZZuQ
XAxb/GY1SXjK2qHL3DWnFeLFYrhxZUZVti1THwjKLMLSKVMAY5CjSJwoNACbFtbj5xNObgOIzq0b
J4XkwONCBpB6Xj/Ks6JrvtjAdkUGvljRc2O2SQqewgzpCqZ6DCT6jFoANxkUYwDEsT/PSn69Tc98
8zSEZ1I8jra1Oukic4/JGjg18bqdWRL7Dhd+82xytMymHIQnGcwEpVe7SLmNnOr8NHYmXVtwv/e1
v1xlb51NOq4GS/mH4Me3BsH+Y+iXZZMBGNExMaKXsU81fe8P0NsFUBWPIWNUmBehLJYjBFhzBeFu
MULYk68qbjUxYdhqvnANllISGzW452irJNBEHZNunVBA3CZl/WqslYSjxXckp0wNm87XFQ1k40qh
JM65vqYN+KT1VVWfjj3YJ7t8RJEn/gRfrCl/DKfZqOVGjRJjUmQG9hm27fenerHv6LJh/UVsYtqA
ALL70g/sKBi+k7dr+q6anHHoiWk1oNuZ/hdqvn3EL1uiAIeiY1B63piWNeXsxU7sPfXmNdp9pn+J
69X7yIt0rQ6cD3k1Akb3lZrD2wGZxbrUtjrXHXE6KxVYPxhvtiP4NW8+L8V/7gvt7tz3lVE/DGut
o/iEFflzFRPEV4eFxSBojh5nk0beSE4cjw0I8SNNW5iEXuJxRN6EAj60ikOnTyMvFVpDXoaXM2pb
b5jmtZMhQpEFbFUYYnJ1PPAMM6at+2cKYgbMm4DoqgSAmPv6wpqcLIQ+0MgP4v9c2vQUG7A/fx+Y
R/x37Dp26vzin4IkVue2GmlkXNWsdceOqY+gXRrGNBPHP7UQ9RqlHi6nYusArk7O6mgJmIk3XZ6J
DGE0aOhwHQmQ2Ck/STaIKB/2695k8hBjOdYXWaumQfPXfNMQS7T6F+66482BK5E8eBY13sYyO/Wm
7CimPt+f+wDibyfWu0gBR52XGtg3TMxLm1NdkCVKGDyyAxV1ingMlUhRZYKJ5XiXc4oCRDp1DgJQ
pSAoK5JIyoxRmfnlLv/XtpuuAbu3WcO0weNxaECMO1ARAu9yfMcpVyzWIXdZoclCcLN8XLFJXWAT
2AuXaYVEhwRU9wElcdrDTAs4VubkfBWbqK9KMW1iH7+ff8LSj44l5YFePBf8SHNwRFibaAzhwrax
XyjevkGNKkQs7aFlvecNgCeWKEgaO7Tulxen5E2jfc0YUlPQrlHwsCjLIAcrGskCWINO08HBVEG0
o/UnPyWG7i1dojpUFRKeeZ879/eq8eyd6lM56Iw6EUoosjxP2C0NphYi3Gj900njac5cp2AtqhzQ
yKhu7hzMu0NBFzNBBLYhvZM6B/RdTLOt4IMPXTopkKKSoH4gvQ9urQN1xxesfl3o/SGclK0wRvsw
6bHyGC33R1Secf1ZOeYccnGeDtDx4sOtF16UkDW499csGzTZDw07TbO5WyhaIk5o0Hd7JeOIxFe6
Xf8Vgr9dS1JVkFlS9/+q7oYI/oJYpF0sF5zUdycdiWxJpT6QKStgAPsgoB79n6YJvZqAyq4CxuCD
kes5CA9fq60kZq/Vdc9Pic4Kc1ZXYHUR59WGZ9s84l4RcVgCudUkDmV/gE0krWiugfK6g1LkYxJ6
OVt97yUrQSlO8ihJgHZ7nLsFISvVYVb1cFv5DgrTxNEAEqn+PGTjwhALs499mcDLsEbKt/kG+E29
h4x3Zmx0d4OQJKmFp1iUFxMSpVDD4S/FqNn5EwFlaMiwN09JdobF9BAq5096LWgVJHfvVY3iop3R
piO0tEoz+7SWXjjdSMfYlWxn4KhKzeWsVwQO0VA+7jJzZxD5SPcY4JSUCNI7VR7IacqET58wxTkC
A5qFPIyuyMXqfy5QLSEAl/55giFPd8FCq9tR+nq7ASs3rAwA4SGBm+TcdTmGU2daofczGs7DA9fi
IM2YZUOzmAwQFEFEFzVcRrezCnaC5qCDG3iAFYymmB8JyBiUUn03NgAKib2nixqtzXzHigfpzlNW
TGCUGG7Qm6UgVtfNy9+nsYftc+J4cBZSZmZgcs+6AQ+dt49Ax7FHxkRPOo6WK27p+pFiiQErF9RZ
abQJFGdnQqL8zp94F+sa/scERotuYAMs4nGUY/NslA6la4rdkZqj/oksRFLeg/Ide6mkDNULTG8f
HADRHif0inmaSEguOov9FmtBdhqDKPAmveDw/zzxo7AvPNErogJVnCDlXinNkQa5nVrOb94Gdl5e
UUSvSIENols08e7z+NDTg+A2t/hyW/0KDl9rRIItQn7XoHsrfhrH3c2AYB9S78wL3mRUYp33nE3A
9tVGn20PLkgtgqZhfSOao/l6kZ6ObWNjh76J8DT1X1l9DX5CfPFhCxpTJI/fRPRu2ccBYnPZvGS0
GOf/xHAjevkWgKgC4DkpaqNnfC2s81y5u6dq0b3lSx6KZfDDJqx/yF1c/H5ebxDrY1JdIkZWZTpt
05uncyMioTG7UUoHejnX9I8oF5S6oL/++ORVntPg2ZhjT9G3HA9DqW8O71ii1JXeGgY4VpsDZUEV
/eA3j5mn7tBB0E2R/kGFItJQRXInSE1pkfdy5n6Y/GwDScdGt+afzf9lTYMi2fhtiW3X7/uH9FiP
apBooQP/IWbB91dMAm3Zqp7e5eR7El4Oir2QyqcbOGX4pw0iCqGaoMxF8HHzBujjAxVk7RUy25cd
wue2Z/aJkKH0l85ZaCJbv5RD1m9P5xmD/m565RkTUASFUsvCe7yU2SYjHvA/IAhHyRJM5cv5TUpR
79QgobCtbOdI56fCo2VoqA4gC8z67Za6PRWzUS40PwZMIpUs/i4Dz2Nk2ieFwtlgcXp9MnCP8HVU
tirdFmS4P9JQ8HXihnFEPx1pDOV+S58MLe0djZQ4tv6AP2E3pkGh8utxthQekmJvktphfV7OOkAs
UCxMGHUL8YaZrrreN776UN8uI9D23F2Y9WJ9CuYAQkBnHmbwYrb3LR+j99iEcBZ8lz41s4s4B0ar
QzWPwtivJJu8CMVVRYVxJ+Xuk6gJH8ugqVxFVxZnX17IvVCez6eaZ0EdJS+lza2pbi/ug8yFU83b
5QQ8xluFFhfxTuWUDmCqIzlEEozPUrjZsD8wYmpRndz8CrcM6vhvr7+/SrzaRHGMiMXgW7yMN2Zg
RJcWPdqiTSBaZhh71+ZzjKZ2I8Y1zVqfItu08xTgzCRKH7CvvePSrfHpmnvWN7BFZk4NInCAZmYU
9KZOM65i8wt+nOgFrQfanGKwp2dOGjs8zGQHGb6hIqTFiidURk7rcToFZAcGUg/lpJF+1N02Wrzm
92JHpmvmpjSv2m7lBYx7epmJTxCEZ1Jj+1b9y1KPhvcpT/7Z6f/gQk2aELubAsFnhGMXNO+iqvBw
6pL0zk6vF1Mkaz1jmIWkVA4FYHzygUamXVvT+r/86ueuXrV7uirZYPxxkwrHrcTfti2mqHxsknPr
YaiH0nfCwQUI6WwJHqLA8QCXxN4yk0ETDg6yyWJ6IUWCW8qVFhdcKSJ9Wxe+5FCYT5Hqat+17dW+
NbW8hQZnqMUsZOQpQrIgn04tYaRtV4B9rsxYvH0H7r+tE+POsmJbfvkRym6EI/TIA36NRzsbk2t/
HOux/y8XydBwlgokQs+G37b+NBEHFEe96+36mQnWJTVNONX7cpW8f1q+UDeTglLKOZoX4c10XJs0
sgsUCV2aKczq9ZtYLKjB2/k/szZMcqhMeYdbyoqet8EmiKnR7s6vvqtIEVqMqPTHijqwYcfGwgpj
8zF/dQSg8RWs1XcOYzafCIpEu1TGh4tahFzxq2OTnMTSYtQvQPrMQBu2tQbAwSzBQCeAQZq1BIis
z6aQZbJ8HW0+TI5CIQNYUArLgpKLFBqQqeK9ixLfsLQm5B8ZIe4pP2pjyfZkMrrT+UgYkzQH/iSv
UoojcO7g5CSECwH/g2TKdc7sf6s1XUkAv4mHATxMTsfNGjXsivVD6JIHJPGVynz2v0DsK8DH2GrN
F5i3NfdfEa0/EOGzJqesEbfz93Y5aWSp2kVOAMnW7R8xmdjnavYfPC0DEYOe24QxxubxJ93CFVV+
ugpmKyO4sg7cwsSRza2JiACf/VmjmaTFeCb3Yf9SOueCAqjgMw+IcpRh1U2m0VGNdK8puKpy2mXJ
m4gHkEXEeRzj1y1Tg+LCLBgZSH8ws34niWBhsu8dquHMfzFf9xwGPCpCnaYDIy2QN9E2kqx3FhHP
Ezmf++7Tq6TvxkDbx+6ebGXu9dWHzWDMTzuZORS+D1gXUw0/NRrfvH/aIJ5M+i17De4ZJZbQdOho
yH5FT90nDl+fcWCIBV3hIoftIGI9weODlDQifchL9r+h5L6nnxVAB/ZcZkzfbUSByzv17eFs6+nW
7d/8BopFp6hOUCorz/z8WppDuTaVXuvgfUiwfz7qEXxc8wAvOsLpezRz5GXNQmzGuKPjwAr1jeto
F2QV1TH63Pk8uibmd5uGhOHypPFidIeHmntxsK7G10jvPFfPPm33YeD/JNrPiN+pKK0w84S/mBBZ
HJq8SdY/1hxEuZDSB5bSPHgoDGjMLh2Hx3AVA42zicNRdDjvBMau4Rkg51ZZDSNeUV2yY6Wdx2Jv
kGL1jPFOxU5F28fRczIyJecCOMoffZGNjYUlaGaE6nwtS1phc0cAf8PAMrG5bFxjlWHj8fStQqWr
A6qMiwK6UZscMYwVkgNH71w1eRv6BZIu5+AHw4oBmEqUXxBKEsX46aKe09AO9HAG9YIA+8wjrn/i
XQuhAhA/CxSX6RptnKNKBquSJ+6PdTAmhg25x5f1PXIy7m9exjcn8SCgx18ec1rf2vNbdeJRyBgR
iydctXCsxqg5DycaJ8d5KIjyedlx0RUaHDkaDbnmKzQS6TccizZMISszzJPJ+5c4CycDkLLgFHZw
s6FywrCx2Tb7sCJwzdBOaJKvS6j5OEFjVXY8ZjEOh+BisRvtDu8wCMqCJfdOHegxkW2AxKPCs5PX
J6/2jsr/yOtXUGP16KPSi7jTB5ybZTo3ofMdRjlvOlkwS40BiFLPiByAydFSIqg7RmvTegZ/6EiG
/Ik7i7T7eozexTt0GF8HwydxEOzu0Rt1QbqOBv+DNX7/bkUwYCNBTsNVCe90yfNugdxGa2HzAFDS
Itpw/2MhvHvhfCIopy63x4JYnbJ5kqsJEeOvLMMygElR6nBrY8Iq7mEpVn03v4cMkXtVoOliaRI1
4EigursZEBZulsaDgqjB5r5m6ms0GtgqmK5ELrMIZ0vUOJHzak97Uanwsv+vyC2gzeDUb5a6hD2H
4Nop1SS3g4hgOzuD61fPlEt9IhsAHCewf2cZxoUjPygVcpO+QywfNtirTGMjRKaPOw/4BZM2/3OJ
YHI2mcBRkhk/OOksEY2Zu1su/kfKz49vJMH00u+FQlnbk2p3OelHEkAyyPO04+yWgAMaKK9tv72Q
4KZF4XLc8TuEq/uWqHfVgcCEcUW7ZraGm8P2B1Wlq0DG++1fmRJk1YV3ZPKpFVIkJUra0nuxxlbT
xMkP6JxNxKN5TbxZJ5hU3jBpldOMYxW1C+CYVGRmeuj521RWaqPdPVL7sfHgLX5HkeT2y4n7YBOs
UR8umIU3JtlzCZyutsuzOAusMZLtpraxiv6miV4NEo4zQ3r8glI2Dv8VE+m/M1JWlljy6TT+Ji+8
2lYYutggqhKklhy7CsOm2+ONDcg6FPeflzWN/qTgJ7shrsB+8dKr5DmZXDGEahE4lbetJRwuUn7Q
0KSOVVPfsuaB1onfhsr/UXL5zCrYGMZlKOcVlYDhs7YqAwLRLnPloMg9jgKv/i4ho5k9eEFq7UG7
39W24+cOH+6ELRST3uK8YMB0J3lOglcNQbSx2TYhz/1TVRtouOGNF6z3UYuuOivy/NO4kI65qr9x
WtGidPf27opOC/i/vKDf8eZQyKdb5W/uxDLY9EyRco7O7a6MiYNzYEuuCzzQt8CIx39H93Nh6xPQ
6/HLd67EJNoht/ILx4EykYCBe1VV2V82upniCi8gNYPv8tdglcSqr7lW7HKYrOSHNv3q3u6zhAv1
nrw7GFTXxnRsKaDQNnKkUkHmlwW5DZ58ke1j9++KM0QSS8BuG/Y4kTzYHNZ8Y/9ftxS8ee5vaYKn
LKUGPANFlrBZMJiitJxE1MM7EcuANO1J/CBxcTlwfK4iU+HHTELL5VCSO8BKoZKfd3N+k2nBGvE6
wyiywjGtU37CJaCKCYLuyhh1PUXjHD2joAkJri1HrMpcpddBvW/N/4NJ/4375h/lHHyQT4zVREdd
Rc+ih/NCcsKEZ9+SybdJe+NbFekK7EkrBHZWwMCg1mz0wmsPzeNMOUnhR3rqftPWzBdHj5vclvZR
oAIPAgPnyZUBFHMXw+gBh5WPxzuwTejYzrndNM+NCSndMcDgjhWIwTcJmiO5kBHFSxR3PJzBYP0O
O0DpbA01SKYLke9QgtO25+gZZWIIn7LdhTBKb9xQZFx7PmNLXSOJz9OUIQAbN7OnajVdE+ntifOy
1y0+EpR8yhmwvgH0qX7FLRzud7Nan6k3wb24jH6x4IOCRIlgpmzLsD3W74rqe5BrciCn3ddAGIaq
K1i8BQMmG3FfNxSZff7p8UkMheW0RuBZjA5UBadfP8nPLZsJNbDFttDx3Y31pg94pH3XV5AsXqZ4
Ul/S2uB+pEfUkc9+tW5f0xtaspSG0XsaOd1SR1Tq4oBqJ+T/Ugg7lH6jQRpktSBTf1g37AbcwYoS
AikceK3Tj5yaOSvX85hQSQIFNIDZvIzZVlwn3lRuV+HpyMas01hcc3D3iuupFftnF6IcXYwCh1qc
2P4rnh9TKsYBSSNUqhggqUADZjS8g4/43hwJjlozQuo9OXEkTrFVtIDy7iAk+711l1FdvP8UDGGK
VNYaO8T8pNvkrW2JXpTa5V7R6JUGO3gSllMvmrQqRkmspxw6+L3ojw1qswc/F/RVO57bgnUisU8P
m6TQ4mg4K9SXbUvywYHtbxI2HWnEF4L402gyTAwESUF1L48sgxsC35nv3ADrv+Js/gUHgr378O9t
L+iwD1zytd3SqM1di7hZRwWDLsBmuPPAnYWRBpJ4Y2c7KuV91YZpkvmj7M3epziJM7xUCPZWsIfV
ccFcDzfTAfYPEaMdr5geyUf7tJ+0UB+JMBDRZ59IvD1z2VW5qRCKltO6YNCjeuiLHJCVJCiF6rnW
eZOKf/elzVM+LS1LlNxc9E0QXx8QPqxIsL2LxlgBKjJpr1xsVv5r3EG7+8YMcHeye0ffW4Pb8lgi
2q3G28tfcikqGbYYnCRVy7oWk51JNawlfPpXvvZluh2xZVkhIHOZ2kye5qLJUliBXtC/LYmKux6D
7cKkDlRKxpG6n7CPG+nFXhkJHK9dhX29uaHGYhziSgvH60/RAJpcj8fBouPr12HCl/UYmgSFZyjz
WdLrQ+KCLY2NlUKZmfc80vnkWuMYdEBJpvDhJu7f0kbxkqTdy8m0+xpHV6Ce249Z57irp09vzaqt
J3aF9V8Ie6DFUOXIje9IdxjEC11yt6kVW8juO6yueknpyQ8neJp30mjSGEXStWcUx3US+tgIgUN2
eiVEb6/8I9v1bERry6vVMBGHNaD2j6Q5PRNOjYPz2eEB/mkkfHuW0EjgbV7opMDoHxwLKU8RD5rs
tRivG2sIiJXDcXchCRDrZCoGP2SdWeahWiMl9UGQd42RyDaYpo+Fh63HERv7RIGkhJ1TVReGaalp
TxxiCJe8G9c0o+Jj11UniFu1j0JQ5jG34KCZcEoQSRH6itEdvtMs2rTDHXZrmKZp+JLv1h9ZO0AQ
iLB8unfCCajPVtu+IQzdQ1fdtsF6YqJj/rU+GZ0+C46js43ah+SDnlbiLvidchjHEmmmei5PEdDp
mn/weVWIgYBFFAvqq2uQarewhnAVvpnulzjXaF9cUUXF3kJkwUYQJMT+TcjRhIQR+zYVTAvaZKc3
77D8aiyVBVYewX3XMStUy4MyORUV85ZoZ3tmIVGtS84lsfuyYQnChm+k/7i7wo/1VQalkOoXj7g3
WVfb0QEJ6Y+hb/0cPNtERn5qzoXg60a2kE/EPiUR/dTa2sSwEeARaPIjmV9ZJyA7dJANPYiNCggs
TZjPoIIRzWqCfAjmMbWaB5+nvahS42cBLu2I2NlTSuaKZqXPYAyCh55FclZnKVmiuEc4titk/CGI
sV3s2Kvg4+cH0ysWmNjJhtyXMTVbRaDmDsYjqBHg82Ay+8UzIsWVM/rZDCUCDcYduZleOPsAWeOx
HOJM/xmNiXpgFkEH1y0dIZ+lcoyXLM9LH7yaxofqFyLfXFS31zW+ZqnkoUTzDmwvgUwQbr42oAwk
mBdUdJCDYUbKEQC+Ydr7TCrzdYStT3YIRJGFAE5NYX9y/M860P7TyRhWNughSipf7lvMFsMS9UHu
qDlGWEhhVxpdtQAUhrug0qO+9kUnrdGJW8pfyXe0vZkmtwwY/HoZOMbB808ki+lZIYy+waIQoiX+
9EhS7MvyZW0hTR2JEFF9JmZnWA9NtuzGFIwafCqt+Mflmt+nZ5v8ffnD34cndI5W/MzMksaH0aKc
LF4cdNDWkMr/jt31rkW77Gm/MuennHfQfNypry2TG+6xWVDofJAd7SnfLREiUuTFdd9d/gLO8SyP
mMA+E7KSuw2xWay2BwBw9nLdfDrjtf7l+Z8l1rOyqj439j0d4DJ5VdG9weUTCFBhzUoJMKYg6H97
Y10mwN+Vvv9nKy8pYlc1xVCzcwvuv0+N/0ZBbRUINSAKS1yj2jGQMzue8QIfEtM5dSD/7tbSTJP5
XTjgoHj1UzaeIao520cpdEixedz7kqXTLEZ8/M6e2l10J4vlUhRxPiH2ASINlnH/umitelLNdjjm
u5+IDpBm/axqgg/EwlwDyzl48H+Yw2WaKFa8GYexDTdcwaFR38EXYxktDK+pSby9gfl6pwyqiIDS
NI+URklEHi7A48eOac5ho3LlXVkMz8yhcz2UPZYuS+Yxc8OqB7S50PUvvJ9BlQIU2SvEcQ4Omd87
+WMZMMxQospupRhzupZzxDZn7IOU0JzerQGXy3kxYyhBnZ3MGVwB/hUF2NTin4GYJ8Fasd1k+B0i
KH1X6z7UBcQ4IUwgVjYTRILLSf+HFzVc1BSpfPQ3yxYcxk1R2vB3iDcVDkcCnSSXKKQzVZEcWrJ/
2X83RUO6nm6eYwlCSLio8cVC3t9HzR2OsDqKZxGzBdSLuSAQ3dOTtjQiHhWcq36JKYpLNnJFuW5E
l3+WOJk2rbkfOOVdQD1erkUJ8MiQJs/48MpCMLZX7mZGKuS1jBdf3IDsi0sHISlw8BVk4AG+CSQW
Y7R+mc5vIuKI9NEV02mHfBW0VGGwTe/DLQeX25GIv1sjhFmAz0Ay6A8QVQzVD2RGVW8ln7ps+ox4
F9tlfop77OtgmcA2A17iUeF44N/x08/JmBQaa9MzijJ9n7xMjcviPyS/n8JNfcPSpreZ4TlHv9IV
vRmG3RnoosQSiUFzavQ3yypCOE+htpAXuqlxi1OguIYfzibcLoS9n1VV7218c73NsI4LtrrT9dcW
3zdNT4+QNy+ysbubWHZU4eomywMx9groaQ6aINWu1GNfSqIzIj4LsRSF60XXL5taucLDIsjXZRqR
iiGvNDcPAeUUV8fqL9BUhVlp88lEKiJ2Yip0FuL450B+tT+O7GZB0xfAtY+epbj+V3WMAyoaj4na
/hBd7MNCvN5atIm0Ruj3gsmbIFWcJLMYtyHx6K2Q5Zu23z9WfL/ZZ4+uNC1hLXoH1t+NGkxbLyyf
X5DJ9LiXSxJoLEtsuNCye/gb7Vbg8yw1VcDTSlTn4kM2khUtqdEClq7Tdoh32h+AMt5n6OEZanxT
BnfaIVti8bx0y75Bvwv4/1kTckQkcF7J713Vv00bxn9WxK8FIIb6Sdpa4YAH9HA8RVnhshBqGo7j
LoioRn3O7wAH9kSiHeOpwIaRdycFQSpCiux4NpFr1XCa1ByQ7TOeax2czO1SJ6Zr1OJIuJtpfa4l
FVFbvU1jZAO7jvTXUiiNyKljNBWb/CQgiYL0FBVVIA63ZQfUevYd24aSawFLzGi+1pI+pYQm0Q36
CcQTfLcCeUZW05dev2Ri+E6EQy6D4H/mTXJg+5ipMZn56o3Du3vQQx7HpFf446k+YHWaFlcbiPkj
sa2/bwJdQurzYbR/CFLygcZawRi1JwbLTE5echcKZycwf0HUePjVSdvDxJP1SGTuF4XB2vsQQX5G
BfbMIi/n4LFMTXh95VZRVDHpflntiSiQnv2WwlssyK1k9gsJIteuzVnb0rINN4etiTn61ShWzi1D
XGJcoPBRd0y7OEkxM1/nQ1ie2lSGbAJGU/76Dyj+JxMbaUmnlA6vEoR4oyThddEYn9kid1wd9q8f
BM0oEAk2jIVhDl97tsP4dHdiVlqIBUaeqWSgVjnskHE6QnWvxGCUItOr9wo6al9e7+V8OUu9cxDQ
D1I6RPbSlAQ3Uvss0R9ATtw4qheMwyDPQRFTN9b6/DJA/53H/7cUTkoLDLXJlrQJnDbiUVB1Cpe2
fauJXqgM0vDcbl9kob3/bG+GeKQltCMi+lG05/+SYchoZwEwRRHFPeRFvISqgwykdyARvBl/W3NM
IlBeI7Rx+C9GHNtMCKzbWPgYqsy9EwicivPGvxLPKMpzXRKvMDbm926O9pS8ebfCxnIuvwwjfqiQ
e0JCFF/PHwpd4aabyVx5MjBFX11tevpw8enEYqN2SzILt//7QJSL9COf5n6aIpUTeDqUHjEFqt05
OFCakJT2wxM7PY/u8MOeUAm8M0vai3726aFbQCfpu4rEIbf1mI7k9HRQ80l0TNqWbIRSaqz+48hu
0/DeVbnDTw5C1OhYeNTGf4Pg342QPs0oea52nS2PjcYP4kASDopaUeEBAu07juOhpM6VWR2HFtGh
x8thdN7dIxSOU1qGNrzBV8+fhise1uuPLhUZ27Sl4pGcUb2OpWCjAh5WlP/4JawvSERIr0G/cwWJ
B+yEpQKDaZvc/0hinWWMlFQrqmekENNz/ZEqelIN1jwFKG53AIfhVSA8XF7tM0S0UYuAFm8C6Wn5
AAumsfF0EKyiCjmMShxzq8jlotnH5T6g5s/gndMGm782Ir/t1nu617qm5c4zB2OED9oBF+hAV4zD
mU2PxefqxmkzKQOS8fR9xFVeQYISB2h/qJhOc7hDGSCAbpxTiQRVz8ovFXMbsoHELrz997nuApRd
KmAyrHWq+i5GWZ8HJYz0mcC2yroQh8Mmd5kcdJvT4VnkhpPDCFDexnPqJJM3O28F3bpPVL+rqC/d
7RBp1ScQITm4ZtcFaaHEpfFkddVae8EfLSbUEhyY6alVpYX9l0NbS0XZ4EIVmUzPX0OkTaMOhbcD
tB4G4AFioEwCfQpYtcRtJpa183Y1/LwQbbsxZTjj4hqmkTen6UXGflBE+X6LMNe0LSPQV/aOgPAH
GshJO/JQWqpFX/gGeKM+YFUlqennRXNegSZQtnXNGmYeRHvUO5YUiXg34/iTyFkF9HzJb+1DW1Wn
HYMW0+Qj+pgkVX+ivRe9tr9BKyBIwurdX/uBckxzRyr9n2E/+FsqkDHhrEx8MPIIXUJJkJUTjwyl
XNzFt9fzs8qrZjYLlAXj6Oo9Qh6TE9y5SNlZbp5os3wOVBDeaEDcanXfqYtrxbkRCcqd51E5FnCq
Aj0FtgYglR47eVsXB9czaEVQCC8PnjZfBU4f/x5YjwZqWh8FdMOh9ZN1WWadwyaeXPUJbDSyB0AN
afyZuyeAzdJBNNZuNVVfdLaVROHDiQNTJj3DJEq70KkZC1K1shl8ZehBIXLyDqCJWB6OGujoFO6q
Veh4VV+FSZzi7HUp5hHc/PmYga49mNLs5uDP177ZkzHjsipMYsZ9/kfaOTIGfJAnSWpXt/3R9AQ/
WNavK501sjMkFOggXWIt9ykZkMMRu+/lGnbs9pyaWmKeL+6l8SExap0t2680fwgRXcPXDm8xvM99
yf9xvpyFZLBg5dFxgGuHjc6Pw35Av0/3Z+FRrwKsNzycT68NxWVRJH8F7M2Db5wXnqlNtHSuhEuC
Ljzu5VzJlVRTyYhUpSSlALhb0qnP1I1cWvajsdDd8WXxlMzlfdoo350ul53UNl5BfTG2ThJlBi6/
BPnhbkN9L9vplK+hOuHOLAnsROnYSESFqGExY+utxfmvef5+vZW6uNPZtGK1fZAro8RgirIQr48g
S9KVp+/5085jT6aUf9bwXOK46f+bBKNkksJhD5B3x0jciyEmKhgLxj/JqjzuWO1047I5BYg5Z0Va
Q15aLrQKt+4zquLgQwuAylSvKEWWTH2EblCs4v/4Nv5iIcBX1vwnTtycjD+sZBEUmXs4hGbiv3RG
fPP1jd8OrMJGxTXk3cGfAy/eSoPNRydabYNRvitHeEvE47l+JXpN5H4Ll488ChLFBODMAlelo6X8
jhP6hTag1u4FKR3cxEBQqN/5bDDrv9PUR+wv378LqDLerBd2SNEATGjRAtA9ulbWUc0hHZEAoqH+
3Rnnpb5BHJ+qMX44N45Fw2Bdk+rpwbT5xUdlWioRLtwyKWjZ9Y2G9Gt6pcdBIQu0NYAyYNp/QREP
hruUe9TngxqQ/xHjaZzGz0Q7rg2DXlxcj3lhddeTxKa89Bdtinmv69ttVaxktDvXVkNKL09TDUM9
V2gmLzGiuIWkEAIs3hw42YL/ya95KQ+VEIh6V+lnyBlwSHm/zUSWNdNYNuJlmVeiOZh9qiYXt9Yr
0eE5ExAGQxUIcSlRfLpS1Cs2cixil0/yuwAIOqQuzceXbDqtH+ybX4erun/8Um6RBjZjx/ipmxyU
aIAqJwk+rIWV+HPCGc0AHRqK0SO43yJBPsdgCvDZ7gFHbWnVd+43w8DyMAdPP2inDiS+geFkyDat
sMujgqafirMltkCoh2TB3wiuF9nMipTsAuz4CfqhyczwQYN89lysJwYrVNC1h22J0ETx6NPJ41sj
dEfFQuB6fJOWOaivje4mRirK3dnTOu46o6gHu14xu6ruSn1XGB+TFfwgya06F2Zmxc2pUz4yLrIF
kGfxE/+bhcRlbqFHB3MVoNifZcU0+KJLXg0tRRNTLvDr5+uMwJglFRU3pPmAY4xyc4hqDiB2P1c2
RK6hRvEo3m3EEi6r6OQDPcWWFqonBJYaMgguJxxvZlu0OdQ7dGWxwAlXzWN3pT8WHbuYeL3yIB3B
Ii4vAtDNa0eToCWn5/QryStN9nYYa9spb4+ZdPUgeDGG/b2PXehW24b9iXc9HJ7UkgfeHYo1lhwt
HEIKitKvjLk5oEPyNDgQe9DceUJjUL0NmplQoWKG0/gIGvF21SV5HXgoK3BycfJ+SG6NamyOjJTZ
ZS7i/rArpv6kqfiQIBOSLr1FkLESy4zis+ZxmSjTjVdK+ySWgzW11sGjoR1BFb/q6y6FNIfn8NBm
evlWvulDSYajGFQw8uAQoa0ELG/ZWq9kpFpIdpXVdlrZubv6yEjK8ODRCSgafuEFs4XtAMaqObnM
EZvHSm1XqU4eTBCnMhgfbZs8QK3CQXSmpAFI7WHQ/iinDYXT+sZAWJo1TXsuxUNasQw7eezd7Lv1
ZaNEHLP77ZKWz34rHO4PdmrXCI6HZBkQfukB0lEVEgTkYkqDE66HJROK6aeryDJmwkUKtDQxUFjV
IHMrNJc4wMqHu64p9Z5geDkuKQAPoDEUAP8GEkukAtMO5g6UzIORNW5ewJasAGRXdj1KZJHvyXIZ
PKghNivzcc0SEEH2kC7sENb+lrPN/Y5+4jPU9vpX6eqvvqo7RPbkCtfmwm3dPgNPtlWjyv4h2riA
1XiLgPNrdIbcjRGUQaBOWAybrnrn+6eY8Amcb8IeGpCPhuW7dDXewDhzgP9hvFG2np+RalqJ47H6
9jf9egMzI50SyQTdtOn5tNx+1RfPNuj6V5RYLh80IfaQuSUG4oEJqKOaizJJ1MXPNfnyB30GybYK
+T02wQ3SukPLMUK0W0XWaufntQ3MofYHMbExU42UV53SoAdXgg/O2uE59vW59GaHaOCeB8Fok+Td
bAhvMqzbm4sp0ieU3HWIWDU/AoDbbNb3DTkHzhHjDvHrTZzYOiqEA3z+E2vQ+UarB0MlwVlhHGLi
O0jfy4QK92A+yHdAJqE6AyXli59MbHUVSXZJvyFX5apg1ExtQCLOZ6apI2QdMsXcUxVUZS196XqM
tF2WFoNbHiyVnfRskRBrF86B5dcj/32IIZDdEqnu68/UQh6O4hxdikCNKgB/2TZmcPSi8hXPzrpU
uNgHuKEYcJ/dxpev7yk7RZUzI791zUr5XeM+mFszaMnVsOJYKrxaPCSkMsuFI5HNsIPobeaB4ezX
S791AeRWkCGnHT4L6aUYvGcIvyJiTD0tT+DNX6ilpucbHCkpK+cEWLzz00ntPBuWk06u37L45T2k
jIA8XvW4whXWYixNKzk/UnwPoEU4qi+frHAu1yILN80cgkXGZq8veV1NfOIfFTbnCOhTDGXfICSi
N2PQUaIqT5ONK7O0oZbiRW9UuPTm7QPE+dSil6Vw+CmzMtMoedTNUVPBC4QK7jEi4EpifvC8WYSa
mcgMCA+bOHAqMHL3PIr5NqgyP39YEqZvu5mausw7FrFrxDq/MFxN0y5sEFtFbLZldOLG1gRFRfhJ
T9pKfvmSeXxhHSU7Dou4DJ0gS/0bXaU45lH30fQm3Miu66xLDkpIc5hUCl80dqkMf4JdBb7ipLok
A02+hTsQeiZKUpok7sUBwDnmCqDnRyTRIa9LBzwo/Zbpaa+uewyM5Y4yN7abgMRlSkJUhGKiftg6
AqfOzDmYQ7R0x/qWKNCZvLr24vsFZPRyFNl5n16Q2vKKyfQ16GqXGSUX7KNrnY9yAibYsx25Q0cw
zw4luevNzvnxSyQ4YmgZ1q50s72LXV+KnrjyLNV8lLHUyP0eePKM/PwR0ugcz5YpSy5fX6ucnk2U
nw+WRMw+kqGFUma94pjmjjSlqGuHlxIn1V+5OSnSvpzTIQElnRrM3CjXO/G1jm3/mRo7mk3+RCpP
3+d1A70sNdGn5WcA45C+J5cm+wAaX3Pq6mvyDXl3eMXsSlqhl9EBywcXQ4C5lrFNhphPg0dGQUIS
PRrJNq1n7AWvQLInQAtdczYNk06AorK0naQK8uCz3RFeYPoppqJnMemxK99kSgj3wYgPUQOe37mF
S9xT+VmBNg6jRGsBitDYhlEQQT2njNEtGboscfVNWHtaf0Dv29IzAz1MqLIxUhwgyldUvBGcdG54
EPtVxdWW0gLCQUNZ+JoFDyKm5nzLJpfZHfm4QjVDG5zWsRBEvJveiKJ90W8Sh42Nmmo7rasnC9Fr
Y1nXYnufpPrYdNqfHCmnAJSwpAype/qDFpH2uxUj++myS5edDTpZdnkMtgaDs+2CQgZbdFG/uEF6
7t/hsO4w0oOm17iV2iZVeKE+ToKBgpGks6KXx5qmdXba9soAQiywVgSILNVFtB16IJFzMfZy8NGO
8/j+qesHkhRlF2GegvERoRP8e/9lgamtn18jgY3S1qVB3lSHJTsL/O4FIlm8kwJpWas8pmE4rEM6
K9elPxXNUzSB/NDElsbnu+Va+g585AcfBEaIkVCjNrqClogb5KpihXixiNnFpMgenZn4Tk68x/WD
eUNA4Ae1zfeuvxsmPDcTql0nAxA82hMVV2NEjzy6NUBf/NoHVs86penM1ntCJd6/QTrR4x0chJbA
70tvGMOu+kqYcK2/3ehRGm15XVdvJakPGOhKHHkfds8ok+m7qx1Uwuw+/wxs9SZsUE+gXT4JvK6S
FWMegI1egCguDqbeh1ULxbhy8noVkKui/3QrGz64VMIMjmALkDQWTqVRrCRGJ2ZID2s7fP1DIIxR
LhYJbDQ2LJ0JTYDPJ/4aEx1LWWCAfpG+5IDBGi5v+PP0SYyLKRbfi+Bfwa0MsOx7Hd0CI8Lmq5nx
JvcFDphH/Y8V9xvffKqFNMMAShWXDWs0cI4R8Bw3ft1Rphpo8Hhvwj+JiaH8cNZxJfxiXF3EeqTO
kS7gFDcEZ+BsfEwh5DnHSrHCDI5/6Wl41GbkXaGKmcNC0Yrktxoy0jjHA+/Fj7ReQlwSD//8/EOQ
EQ+tRjW3RsbHOMxAxjhmWj8GRFR71/g/e4nF3z4V2bChWjaDWcrrNmAAGaOxmKIEcufF+d7DimLa
kF+JzWGX7Y7VeAUlJXpYv23y5XVbyw3DPZNI50LZ2mSVWFI5kgvgboxA8PWteKCaXlYe70yJsGRr
moRl0k5FJ3PtmmPV4wF8PEiCXQZFDJ7S/OoxiNyH27V53JRpQkqSCMCFCu560mAUPISFjuRhZqPJ
+kB2bK47KUmD2m8lHvVUIaPBhTiti21ANEYLQ3RvVpO/ynk6wwCD0nWhmyDcqXwQdkC1qAvuRl/+
K1f1hopeFaEfdGH1Dh7FqpDkUP7k7C4JW/hx9/U5OBRg6o0Dp8pgy/+vwJjJ/V/VcrUj6sKGKNlT
jPZRPewrn7q/LFHwQOvhwAu8tJkoQQmZsWawWcsbfp8pcrhnG7Qc4cbQZ6II37zc2t4Lrhv/QUY4
SGA+eWYyfCrRsc1JPHPi4N6OuxtFh9ywy3rC5igvXYGjN6kHAr+ipLI9Mo3nb02egfaFfq3uWteY
7BtvFYvc0CRAjpqLs1zkqPvRKp4yguABzLcY8BdaKoRg1gypHob3trj06JG45zDM3NL+Uq/FTPat
hNMCTBAwyJA6d9H1j36LnEE6qOlOew7vjowB2gyRq2ZSycWdAqJn3MOugn1n9xSAqy6MJWnsue7p
xSX9fAV+Q/leW4oH4sR25mYcoxJeJXNiUt40TZkNb37f/2omu7Z7mLh1PggzMvDxGWycVNYtmACG
HhJEGuvbmy29sSiAJKceUeWZe3O6zPyqnlKtyKKRaZEis4mHGZCpskm195kPY2sLj193Dn0Y1mJ0
SpGnCCGqH4hY3uOhb40lBA5+5bpfKYmo2kf4QVmpAj4c640mxNjVTR9qT4uGom37cEdy8q2KCX4p
qSucHn1169olaaUrX8DU0L4QWMkfIFXiYIEqt7G3BIw8O14xVJlFfcEOscfD4nXoIvsaop9ARTMv
ewjoOLw/uPYTXSt/FXLIELNHaGKcDWcD4qY9jp3jgZwm/1LN50igbLHalj2sQiVr3fgv1XpXvuEC
psGykhMxrBvsI3lqgveb6AsMiCCbIMhr8Vs6FHP2X+q7YFO7tXRqAIal2ZpAhDTQB92Wtlc3WZey
eGeXNytp9NpfO6CtUKOWiHDCUSExiZ5kQ+JEeOkSQB2inzlnblrxYNo00NljqZJph3c2H5Y/mJPJ
a0PhrboF4kkoAKIqqpPK8MMiw0ZZvIlzS+iUTP7c5eA8OjTHDHG5r3qnklIfWqOEA7/kg3hLyy4M
Z/QUJFGMm/0zUylSk1z7oMfUjVORfqGJQLkeKcWf8JD8vFSwkN0Jv6mOEeHpwWhO5UtiiO4DSJwK
TjdXJU/MNfN+sP54oRogfNK9Px4+9L8BjG5Czm/eFZ8DbGyovRtLgaHy7vzbiXMz/USHCiAv77hW
5BdToI/6T1+Aj+o20hAoVXptN2KyIaTU1PqtXSRZwHjEdvO68Z3xhmPBNnrv4bndygalXeaUn2hv
8z8t0NpDeHxdH99zAJ7AUNBgN9uut9ZeHS+0wBqfeEkQwTyZHWBkCZMSvFeSea2awuR6rGuSacv4
n9Z9dOsPlDps50vdmbm88OOI6+2JzTA5F4W8SyeWgF+92kJ37dmSbQ8KaK9xxsQQUczDhwgN7J/P
C1jggxu3j2SAO+ZeFAKIefOl7p+w3WG6tTBUPgkjlVXlxiRn3zBOpT2qq6wgZdKvDeSowRn4LjrX
l/V7WKptQrCaWG65B2MNycPWdohphMKEYyC0OMisyXcWjgVfOx3Y5BJpIY/MBYXU54h/ca0AVeqs
71v2tbdNSR2tUI3BI43rwVaAxIR35ysOF8Zb3ypgvEygBZlvvYqukUfennVyIybVwMLmLBpOgusY
TywOXqs9/icdGkrBTKxGwz6DNBaJyBa5RTtCXFRyJ3/wywfPOm2mklV2rzS2Cl+uSXyEezYti9my
kN3nizyTCveX7//Q//uoglCwl4pXCBYDllDaP41aKjFUku+GNtMbFUzqIi6t2wANxLuwKgDC8beu
/vRSpW2qucycYhSaf8Ik4o7kB4Rs71Hq8oxdQBAmoO4RPyuEUsIW1K/y6q8gtugMya7k4xCc6JE0
kMQ6eY0Czxd8xHzCO10lCs6GwnMYN41XPxwcBG/lqDQ6wx+8129fH0sx4ez5qNF2/qn/qSfjYwMn
23f3EBAcfI/4iEXyvFrh5rIqSxBClvkEPmyFq0kKqYNsDkUfobCd7YUBDO+9wAZ2Txa4McDU4Y7E
yRNbqmAchh7u6F989pnKSVx2mr/8d4ydCrFP6kYxAA+7Lk4mSjC+5liFbvTkDaYS6HIAkhm4X40/
PjuS8yyk9smz9RlyYtc0FseGsgQOLWDhblNi1UAZ7k8dC2QM78neSE+wajyuiDuJylxe/vAL6n/U
WxyLgRBo6YmvwCq9egY4dTNAlHr1j6K9fgdAlXgL0WoUsBxnZbgG/K/QDywazuN/BzmPsc5wOAhP
hKRZ/tMC6ft8jl1xhJl6eY7crdsy7NCb4W0LIL3nCsXeehasS5Hlr6anj+gMfpYJowbxg37703Eb
oFKv4nc3UKlIW/Eiz9JUgyJJ6fEQ+JMKWya5+RQEbC1zAzyI6yFoVkqKxalEnn7+cKoQvRMixR9L
oODB0ulcHtgD99NoFr8rOaQ0U6uyUTlYQjl6umdFMRY7pnBZTncxR00xcWP7g+TgMIc1gSZX17n+
yhJmPefL5h2g/zSfJP2eUxGEelZbUl0IrkfkaBQh1+CdBwvSmP1B/m/DUolVgeGnLHWjSruzZW1+
znZP+0S4FrLu+PgPIcufelyihB9WUdUQgiohoJ0ozX+IOMPP2x1h3wDscjOpXqWEaj7FbuOOW0e5
NC0AufNHm5aJO3Lk6ME0ACn0vHW+MlH5uThiy8dk+2+J6iXCHE1Eeff+mxxOj0iK4Z66p4lDFret
sdfPONPl2Y6g/4TXGyllBxZt5XJ/WR9Q8azboEDC7MruHBKSAr7gv3S76GIB1ydWPFhahXLTehAV
YjuI+6OvJhi3Xck8ovMEOGL8jdFMfdc1aGjXtBBaAoJ2p7vdaX5d9kzBf9htaaMre/FNL3Qm5V16
FHGRxzUXJYQa55nJ5wRkWJ49gmlST+S3uJra7CFTKIAgPNeyp1yZfe5g/d1JT70FQgS7jVMW18No
xYlT1KyAXyoMKQjT9u9I7ySGN1gl+29Vq0bsbtmAO6HpGYzEhiZOO17RMqOFtzq2GCgt2LkyDIll
yv1zzuqQCyvsx6MfygJCpTbdpQAYbybOPcXQMTJ8VN6uL5IIRtKb3QJmOT24H479lPb5Vw9gaM47
bczswjZjBMtEE97rBUMM8Kw7NUzHpqMMB2cO24Qi8lMQofdKkB2FYGkX+IZ+A06vspn3i+vqCI+o
iTij/ZRoiSu17net6czQ3OpXdkM1QIYVI/BNk5cLrS89JY+Qo7jS/g9seZ12BELhlql+zUQXb5hh
NKU0cawfJNey3DT6notPmhs2Qaf/en5SkMZrpl0sXsyAtyH1FKf+N4paYzmeWRQfDl/EjvjTNh85
zeTXr+fccclPC5UHAad5t9UtqYtXOw7Y1KqOw3/1u2AyS6IKQB6IMVTYkPzTN9Lj2V+lB29Mzdvn
5XZy77iKMace7+uCmwq+GXUK7FVmqzX/JbjGdBvQUVV0kM/9XImSlk9pIDis7vzL7S3Omf9K4OL4
f7GQ09a4VDJpN8LcHi8HUFcMSBYp/FQw1goba+FJ3bzKq85Ls4GU8YPWjeq+yuK5cSvAQWcvrxnV
4fIDMGzaoEcJ2tIZdJdXaQP9qa7oFvsDrZrgzYG66pEKFb1+E6lHPMP2QpbFZYvhjcq3Zf4srS1N
XCoWmtYLs3WG71wC4mNLVrZHuCbPWCNFYYYkjzEyl1Ay97m8EmZ0m+rMpgpU8PoX07/9HfpHjwcB
63F12rP11k/pfUiKEYs/MczOqejlDV+xsd3BTpxorb+muAdw37XbX51SM+nDbtenSRlMhNzKtMAw
Jp7EBUHcMDLnJqiLPW+ZawIe/mcHNTBlqhk2VWjcsLRkvUam4/IzyQlp5wBMbwFH8p2ZiaUOPXDa
iI4AH/Zc+JFTRVeKPMEgPY47uQzw0euRLBwm5lffqDw+wDx7COao7EOqIQZF1wmKzMQdT7n+IXVl
NNERer7d4j4Eb9vzh87q3NX7oQMS2cZrG7TF0UOYh/+/gp+jBBWvZ8kJbzc6+d2iEMTaUi881hRu
v41JruC30U94qchuqib/P+LU/WgEmJDCR+LPuXeaihyx2cj497azv5m6Z7jjl70NIgqHCr0eHwtI
/v4SS/z6fqfSRPD+kVPH7UgQRlISZHiDLwyXHdt6494t5N3ZqTQUsUq7YdQMtxxqbggCRvdVz7NV
XHXVBARUT9WV6P1PoN71t5Os6DyatgrZ6C9a7tenlz43A4KW9eSIjr6OFUgTWnKYhAOLqxNSFPKb
p048anzgFEXkoVrk/wQpN9vQxTp9zU7zM/5bPwLbe4UYIrG18wXIgs6RYienSNi8AEsRXlN/W/vE
Us3uR+iH9ch3NExqODSBkt50n1F+MSPr9uMrMVLXmcb4um/87NTe/WMBndg+Skvq4ZPmNWdSIuPg
MeDbmRJ2DgkjZOWJrdXnKu2f/PKU4f/FKebz/SjsNOLfSy/Acy4dFcf4FUcKAh2h5JFME3BihPNe
95XM3rMvHkfwxCxhljuVNGMrUaEJrqcNovTK5UYL4Cs9oBC7W0xnE/yUWTL/qLpLIHYezbwE6QGU
56zJEGR9VX082KVFV5umeMkM/ZrT8Dzvt+2ikDbzgrAvQkh1yQfu/xYEIyv3Y8sOSi4Etz4lsVKP
nT16eUhOlMLKYH19CJy7t4APFFSPRSQNvk7hyn96Au1pu9E8+e+uRCITnU3fe9Oq6IZfWbgvsekh
9mt0BA6+F5+eLRo/Z4COTieCYHh30w25gaCoGJDr2iKa5uwlp1GpkezLo4e+pGp8mjm7xM9J8W7z
f78VnNKV8fObPMTBIyHAT9cv1gSrJwTqSuBbzDgIO82kC7K0tzCf3d3HdiiyV8tulEKNEYDaDcLa
R7zX+gRDteAzwOrI8QiQMPDUuV0DT7bFFUnSQ35YC/XosW4pmyfFYR7msefqSr1n/qQUoNRizvyA
kZlyJSbvuDZfvcAnkirqfGyt5dPTi0NtB9JI0UceU4VARhbo1JBHwxAKr/zGOu7w8FIKHeUfBmAG
r1Nvf6Zq1pUlc4HtaBgzGVXj7mLDcHwLqDXoV0edQvkYidUL0XX5pOW6NS62yoE2nLNpj9YZIYeE
pvs+5Lgp/L3jC0D5PIGFDRpuyb4QHHLuOibwWCEl50fhmdNo4oWNMg5SlBHTyvpbLosLMcyVE+61
F+4Rz4u1HKmIN5fi6M3QO9L7pAQ//yIvT1AF4RtIikj/eZmooKhyRaX/4DdcCpPV1JY7w3YFzDsT
v1aoM9leRRMDLqF2U2vCAVvrzZqFGDvpXJOKLodio7laWxgNmGRJyg+jdiiItYY2kpOU//zAm4JW
cjI3L0pJssHwkTdpLt/pREIuTPVZTGHCN2lRNPdY3aac5kT73sdqUIbLodTyPvw2iOkEIdPhx+L+
zYJbGjWiflJzvLUaIOwuH8O+eYTOVRwvSg/WSj97h90CdC7N38BSGMEkS7RKP4Wbrnz9Q5AsXQxR
TB6OsnHxifNolRgWJeLYoNeHA16roZmMjmUPZIFrSFVxGBjKouhbHgn5ztL/HikNLrz4xa4xhaXs
Kw857kOFwSCNFfbfCA3ce7nFULqSSLguXnHTG29RS0esX//6ND8wTz3/jV+ryJVMW/pJxUAdmhcT
dQ5yLRmKY2dVoYCulPgD+7T/wEVw9sQoCYovIZVUjWY1VuDjtIxgqdEeqL8ObwIJzNMfCRAI6v7j
xvSdzDgWPItkEld1kUpee1pYEIAwry9reortCXNOTp2SPFX3aaiCSyChaWMrrKH89xFw0hUgvHuw
O3RJW+MGnTuVFWzLLbfZNVzYHcyOd2CQyn+hM2thfkB+V53pnfJzEK8nNT0FG1lrxs1wqjkiXpiK
ZSOQl9IGQ3mi0SoM5oO5wzjs1kFulIvZ7jHq3rQKr533joTzTzRBGM11AGGPDSzWCzS4VFSQPPbR
ZB86Wv1c9GQBvpustcqOlJkfwE/Ck2tA9m1vK8G5dAxTCMpOrKNSc+tazOAn8gD60SFHLwt8mv4m
TgyNfODMMt+D92xaX75uSx71iN6DpiLXcRqiobW1aLuDAk8wrv4gn+fbwC3GwWZQ/Skpx6K3Cexc
OHlbaQpodyRZE8ijK+POIzNXWVuHV+HJhtx7Vf/D00nV/wvoaYwVYQKjv3NBLaW4WSeC/bFkvXro
Zax/2HlyyC/YdeTdNA5MRl/9bTERnO2mt5B6b7MGzpmVLwInStnTJKKJXfCeIl3wSHeXbdUlS4KF
mWEDDOPnwEcYRZECLpFVaopPzBjrmPJB8Lye26dAv8kRcoR0Akiho6bNmPu1gXiDhgQq8lk69gvK
08w/BK04oaZ/s+lz56VcXcQCDGrL/S5nYJcxss+HbsM1/FyptgJK+Oo2U5pYpN/810b8rjNftSz1
CQoRFQAxnzFQZX4ikrZ0ntdCwke48h7t/S1H8E1Yz6YqUOv73S25/1ecwRl9/OH7wEZvBlyMFgQS
YVRs1ICwt+/FRmg/VryHsgFpgxts8XO0JxEcKNhJB/O4HZHbpAMILGNhCV5bUh+2E3eK68GEdwy+
vh+ISMf6nAInZiZld7LObZwT+XQxAwtRvepqSfU4jSilEfC3zYW/twt6fwkpsLUQQ/T+/0r0/jwU
Vb5X8zPMz5WY7Zr2/tm0MPnKtv0uxz+8o1sW3Q75nj1kNrxlPh7Xx5nFAMVuIqtPLBG7dHwAnTW1
s2TxijeBIGV2tzYzHHDCQIgd77KveN40csp7NA1+43rmE0MAxFKIn1WITgu8Q8bu3y8Gdl/f34t6
hi7ZrlMTHfafTwEeWWKbDqm2yWiZjFUcNv6a9roZk18Mg36SkwuEqUrRw7lQ6/WR5CQq0OCbKuXO
omtyu1OrKWRYNVBiemvRxlSR3n7b4iRASyA74TYBfxPQfITEjauucmcfkgqlxa2kv4XJ74V1bg2Z
/Qt6rQo+KnLziQDHgiIes3v9khJlgeaNOCjP716I6Ov/M3my0swW4Ti8N2J4UXdW5JqsaCoVXnha
R3kCaWrFLCSizF+BOxgwcjtaO/Gnm6uEueNkkb2u5i8UPjDLh9lcR5RMnuG1cIOYgiv+0fc4eyWv
NHImIpZs7fcY0rmGgYlVfaDV59CLsmxPrn/85EOWxyj90CYDL1mBVoskhXwJramwQp+AB7SPIdsU
3s8NErjjm45wNk1kodGKitQJK0F8+DrjhTZnCX0WdoD8kokMwvDfZ6JNSCxpuWxH2XIfSe6c8KiL
VJ3G6xvCdRPsvCWnN7YwmNQZORl1yPcx2bhnJyyNDK3wYKeRlBXiMj8de3qPnYbzcDpNidNFSTly
C+17SuwGYTMb5n7H38jXzjPyvkqSsqEH920LMqAx8LnX4PcQXg0XCEn+6GRYAw+kaIA1Wg9xFgBz
aRxo1gEyYcd+Ti7quVj1EkGgblhKQoeRg3wvoB8MRYqy6fWw6/0oEcwo0FDGkdfS67Dr6GkJJjj/
XvIdYwGioDpmjO2IceGODV+L3WKDSoXfmcPuJkDqraTwFoFWs0ID58jFD2hhMCh9nxHUoKwU7BaG
thDiJ3vPWEO+UaZbbWAXLl3Enid3lvvMCoMa+Loy0iKRwiSw8iR/U0r2sWDT/0BL9ND4OWkW9FZq
qGPhrUDf+2nJPssRDEM2fUpIfQ8GT36J5xpvOZNzZkgXhdT5+AVuPGQyuyZsXHHmMSIJ1pckYIiS
NgeAv+1cPRb3n2DbI815L36eD9WrvEaCTuZz1fHxC1fdjrvN6NXGGTPNGo4RmwLUBVlEvHeyUgg9
ZFXQtZZHJjWxPrr9hhd4U7bLga7jl4fiIW566j6gWGY/tDrn131eglmHLyiH0Gu3TUaMkbTml2kv
H8EkJlg+yyjjeEW9GIkcE7r2df55PkvEZOsAJT9u6fP9zBCz8WWswBeyWIMBiBSyL9QGuS8AkAmP
roXZkLwuEobVBDOvUeC0WgX8D7fNrG0byLK9tLAdKeo+xF3KHC8p8gIwHfNGQfXP2dShZONUxpQv
3lN2FBITJs7wavYN/0ZTPqJdo3JbTHGy6iRtUrK1cwPaGd36kYvBDPFAX+nCXwrqnRBe3+jlp3wM
StBfDCbXyIRTLLrVMHSoorCPONs63euvpAwJazSobLPqQzj/ryW0HnJxK0lZtFX9+Ixd+vPOeM7Y
czCX7zwT6eczAyW2WJUdtEZUZoSx4rW3VyzPHTlfcZfMPd9amOlzOcKMt0dGAWTntByUHkqQshue
7iy7+gtdYmElI0Ksb40+W47AsQS73LApMNaZzIu7HMCqLL0guOFqO1fC1vNp2rItjIwEW8LAoace
BnD8vJBt9dRmHYKlL8z5+ZS4lLlJzMdAot1zPRetZXDEjmSRt22YfI4nXsXZdpQJsBYJDcZ/sdGG
vvkcgWVZT3/097Uk/rxNtIoXm7JW0YjY1nCLCWIkeVtLe/DK7Taq+2P/4JVfAe/sW7bBRxz6XyqQ
1fQcGzE0nCmqhFWp00hgGp2nzKf0PMcVsBJi1jtTx0nn4fqGGIK2TCN2NxCjZX+w5rz2H33/MpwU
8eHa48v6lRhm5iBOEKR5XX01NGJX9Wu+sHoNFE3/V9eKw7X1Yz/WbkL+7yRsL0YJvHHePnmV9KHo
9yoPOQlUbSXnJsfst3H8gD6L7+eIKwUHaknDas5LSTbdYsS1MrXfSNv10AaGY74kDqYDGKu/rv9J
2Xq+CTwbfKV6iddayq96hMkekemwP5JzEybNi/gtEeWZ8lysaUDmtztZpbX+z0ewjCT+Gyp+v/eT
ttgO+6Xit+Rfaj/2//OlS1OgVMxKDvD3+BtL7jcjMkrJ/k109nuc6tEWZqJhocMTUfbu5OYCPanZ
V8woMbn5IhY576AKCEwTWstyFhsudi1yiHeg3wdYoYiov8bBEICFh8I56uhELLRdFS1cFP6bWzqw
zkkrJ1ai1EMRNrMGk4hCJME2xMC8wP4BMwXFAPtQtt5VhR23VoGspz8QtTF0Zq70C5Aw5oEt3Cad
ktzLWPUVUpku5ltMpT0ntgvQaAWwgq8uT2UsfkW+vblnowoEIMOFBWVwl53HD5XeEMSP8uxYjjcj
fESD/7H3rcM5Fw1T8GRJt5IDmzwXpjfiVFHFnOe4E3nx3XukipGhA5dopYokgmM6aPnD/4nv8KRG
qR+kIZ666ttBLPeW8ed9lSmeYmAvzZ0OD4Qps57Fh7ZLYWrXFCNCX14DCChaiRV5+DCtphSFKI8b
Ogz8FDhv2Ha7sSUcq4TXasVQT9T5CNLFEtgIXSjku3ONeLqt9eV7+6quqAOPAp8fy83W21yW45qe
7JzQVj5/6pK2ld+qc4T25zGNPu9olErqlVRhOUgnLmubFx2jf9puaF3FgzeSIBsWpNHFyCddaWCD
soPCnWfam8gx+GZtKUkJL0pzAoy0HAdPOhh7nAkkn01c9b94dnsOFszzPkxE3SdjMX1cufKkHuPg
OJDO7riU+p7+sHvcFZIRe8chX6otlWKuQi7vSt2wpmGf4TfMbkTIZSMVzS7QRVXBztPqpP/5QVRd
qbuVllO5H/j+GfIqiGoDVgueCxA2lzBoQw7+hJ0E9Ewp7Ha/25SU8pV/44rdoPFc51Dxgl9hC+la
YowVckqFMERsWGaD/hQ8tEejlHdh1dVln2SmoC0Vfl+wPrCuvaRwPDWTQ+F+X+JJjgWpVIwXZRh9
HF2fFThVbrE0Njyom/mQ/5lGygF+9pQuRE/9bWNRIaqLPz0gmERzbwnqnPUVtuOIcgctKudG/Ycf
UjHgOILPPs8gIKq1oWpw0lwRWmPjwMvtOs8yezSdybJCvcrEQ42Yb9VDnbp/0Xt3TzazY12G+Vwl
vnsSgUFOl9p1fwjpy0LbmRJn20UOB6jv0y5JL5KcrZg0OBzm3bnAbe5sLpQGTv5+uD3dB41Q6YQL
oWhr1maI47m2DuA31nit0irg7lWnQHg2Cnhhm5Trv304G+9osLTWqYtd/TS7EzHG7B5e9xKjNDFT
jXY/htGfrMAoD4WbjQLCbTFnFfL6+pPOu5+EPQ7MGpD5ywHKRJz5cOWE7zHsSrG7OeSZE2P+BSxA
aN/IZGHDnx3y+rkThDlZyXfidNJhlnkOKhq2z7wRqMh0bAEFOEIZ0wzvBfWVUc1Eii5Ys2YaOKMn
2x1NE5Zh/6hf0Ds/udeRZJ6v8runksz/NsRsELU+X25PAWerkUmaDHvow+9FewJylioHyoOflbC2
7SOOlC7UR3yz9OCMU8Ei2SKWmh8p4Pu+z1zZwzO8x6oQVe1XOgglCevLaiv2syi8tc2POVZqutO8
CJRV9N7/MlpiZlHdWxIWsa9CIriIVL3HkwJMNt62XksyCJKLDtmPkR3sOF7f3sZBpJVCdDi8mW5u
9dyMkffnYCUAl2Kda1fB8NMrWOfSJ/ZbRQ65yDBVlwT/Ctz7bn+gvbzOO1CWtxXNIq6ma6HKUdNl
0v0ek6crIQbhjTzyr64FcCYIGyFk7MoCou0gKNSZybbI7Z3lyHBsVmUTzl1cevnSd47ssXiJsgzr
ZD8HPMKQt032T9tT7ZGBNXQs3qVn/IX5HRaD49O0W7fSW7F0VSPtmfKqZVASA3SJtJ/VYtNdflve
NntvvyK5xqHP1eF/9O4mPORF5c1yEq84/+Bgfnk60O+fYT5IpVC+5osGEtq/Ufa2Hkybv89IuPZN
gVHwrxPTP34binWABI8U+dd5SrFjdq4UXMvbwoRQD/SECTxipMQ7Rwr8uqlu9zoEUcgeC0esvoH5
IdppwXHlCE/D/KR96nPRxaa1QT9WSB+FR2jSmzNv97yI39UU/1jxb6fwL520sProYp3ovH0MnfnD
aTnFdsEQxX+UQbQeXJGobDHyNQ5JiS+2HaiFbmTcuXDXbVJylrR1NWYtCI/7j1khQbMY6PWr16gV
jg5XUuY/DWCgkdI3T+FUxDDz4XYD67BynoLB5Kg8cx6G7xad8LkK4L8ImKB4DfQ700hR/jdOAV/M
KsmZjQsjnrmOUr+1cugU4UE8+2vRWK0ulxA/RPM2dMgSEyplwXEiC4qXI9p0LAq1sliQWz/N8f9Y
3YPkzmq80y53ma/SxFzWXZ9OuMEem5ETlLDuVgVpk4ed/8+CGp65tGWVza1nz5pHT5m0jCd2fPlK
0Wf6Wq3/VbpKkp46KBYeVcquoZ3TF57P4RfPL1rmZdFguuUSaY5ZLi85jU+iI91KDQ7UW2O9k3+Q
x5dINtHh1BehttRIdisUGnEpRC6vg/H5yIaPn1QmqRJEyFdIEEy79euBKRNUyA/jJ+39x9ocMO7c
QZEp6Hq98kRCAtJXXaVEJpeb2JHsZmUFv3B08ANvRoN+ZHfmPA299/IF2N/0mmRj/WTnneU/h/AY
FFMbG8AGZ5cAw74QPu6B6ksVM7FB+z7g8705GAvtLGRHlB8FjceBZ7Z+2f/oHDsWPIfDcZgtpuAg
CyhvIhspFfdKY/OZh93lO3Puwz6OeUeO9ChShGRJ26GZvTKp7AUxq3D+sIyVA6HaYf4Hpvjdmr1h
PER8nhkdAqA6FLOzsm5y301jsYPwTKnB+yhLIL+uHLkfA6MNRzhbw6zfnhGOAITu0vGs7RvS7Tit
Y6NbglMKGlhkHL8rBE4+ZcB0n2zfQIxwi4sVjSDg/aT9K2eA9avFc8m0wJ15ZsY5LJO41Y04C3NQ
LhPXoge69j6OCA3pXmE5tT4DkqdC3Bm6JXfkzMxAjqN9QGPdRoKoyvMusCijS1qJoy6NbFumSV7X
tIDoS6QL/zv3wcoSB+TiXSlKUiqqJ0XxtoBRjsTsdaOKYUncqAiuqeZ3OqtODCKOdpmjnnvkbqr/
0Q21CknioaPR387scuhnKfq+npNGwowu7tANqFwTjDpYBr/rhbSzu5kA0GMckuIb1oZmIswxCPRf
JIWoYhOvn7r8vIYdrQCS5es9cxkAlHjTUq3lc8/LjCynepyPPCUOMU4IEI0o6rtG+q4CyM2Rg9It
vLWRBVFjG0ncl5tpDUEQwJMMjO3c5gSUmYlAJjcPfvoeV8YCmsiH6y7nWNpcmb5342UKDaMQ48YX
LHWlkU3ZVSxd1Mzxc19eId8MDSFyd+28aWLhO00/4VB4tu3fBHUI5phHcwBQZDRzSeGbtmt2TDvr
ZhtIZHYWJKzvRv4pFcXBKlByGG3s5nRGTNokSce1M70MViaEnNoxv2T4mY/CF2efM5S0jcB2LpVv
P8GSCbZ2ZTx33H873dlbTVk/lv3IAVL5ublllPv/P+eXhkhMd4z7qyS5YfZDkxZ28C4tC9+eAgLO
ulgPAtVNXmxF7k5oB0rmt/x0kDS/74DRo5XSHbQFqHui7z5L8Y6VdP+flzA6Vy7j32Sq60NG5UFu
KVXg/Dd6BBVDZMYhnH5J5CdYZBZDemsFMaIVBuIJp0abRKaHvNCZm4Rm0cD/4jRMXt0SFSqtk2PP
fcR41hA37XxfUgGxiBXWHW2CJ7odObf05ZsyocZ6meA11lsUhIUx9mf2IV4p+jaJPMDrJNCHx1Mz
Q9i90eO8wSOHiFtwpROdrWN8PdGG3KF1CjY5NoNv5Ddbf5UYDyc7ZPIUgqMJmGnq/Zfbe3uN0bZJ
IH6u7tQu5OmBrtGTzRfkJAmB5v9FPWsaZBhBepRrxFcfuvO9MN7plDDqNyTW6XZCiodt7QHrFivK
wxyAzhIplamr1rUm2+iDbCLuM0w+LiLjt+Rc2vHU98FqEQGWdUxzjvtzn3fm7D1R5sCUrlEcgFm4
l93usXV1guMoHfVGSu2frsaC3EnGG63nbIQ6nNgNp8Lwl4lDLlzuYOHit3z9hYLMVIqVLVHjn3CO
G71LpidJqChpugMtsrA4FrPKWT5tP7dAmiVtceOlgJwCwnkU0srMX8CkbiMh7v8h8VjYFBNu2uAq
TNXlg0pA3CBrUE15df0jom8LtpctMqfXQGFUeTEAYDXoPiUmV/GJMfN7poUa/XUq3iMA4LfSp8PH
b4BgVuBeCl+emenfhdYdVLD9UjWn9Nfzai5ENha4W7Pm42gPfYqpdVF6F3QuXbuF3idkJ0WbBUpM
qGEtnnz71xWrMv3z5y4Ym+jgLxdHLQPpAmINInv4M2hjjykMvTQyE9cjaJzKFji/j60y/iHJIAZd
5z8sbdHq616DuwbcaNX6+OVW0gTwBMT0qYEDJ2W8Z+tjff9DlcaKZ7oRUN4FdG57XkRYc8vvlUuV
WgXwadBla610tCBzfeavWYatoYy8fnP3X0vYkoABtsHlwk0nN5NXombZ1goAgoQlfoul4B0w5Y5E
Dni2/K8uquDg0um0Wkdft+MpejPyCa+5iD1ZgdjGWht+nD0l+TAe4tKGj5GZfus7TZvd7X/GRlnk
ImamZcrXSh8Ri+A5vOL+6hyt2DzaJX6iuRcIa4Uz4gAHbdHOaXo3KmrF359M9kKDCC0tMj3zLndH
KYYVus+5n9hwSLwAkosvb3Azi9U7YpakDt3B7xZ87rrEEIaqNbintcoNDU0J261pL51tW0iAajZF
tEU+t/4YoDHymu5ELup4fndIE58TnorpkNlJei4ZUGZOGekv/5NOY371/4EvqfOsMhJPqZybERCe
rIESy8VMOqDe8wcu3s34LGWwvSC6Fii+CHYvhthFxANVONmht5c7PZ064Pq2fKa0w2F7qRdlHTQZ
czIbj8MRc26l7Us1MCHJkflQFBDZ+roJ2KmRRtNLPEAJHuAcoo6PkzQFBqvLfBjxwpAjUqp5z6PF
lX5Pr4rBcdNboVJDckdBUqpWt0QEPu2HtKx8fiULTKbUYy7BYEBZsIsWk5RfSISGbIwWmPMRPB3m
5OAipdF6Zk8zYNbi979CF/snvpCABhhWNDn0EzZw3OKDVbP3/fpCGNSr6JFnoSQYyuMG1wDsg3cF
KZYDz7Xt/GekmJFa8sqWVqDpRELfjVsYsFYKBxIGWrEOVIO8pPGretEkOn++4xPWNyhURxYAMPVE
YJdv0STyujrqVEpciYjIV6rfI2LzMJ7+nFN5c/G9qlgW0dt1iWT+7pAGRCtL2mcAsUVglFlvfhAf
2/e8UOahEiwog7/K7hb0MzQ1uW/XY1VUPGS27e/ml7cUUQrI+z86f3dZsqTlO8fHBSadU92ImPHi
mEqB/bOnU54nsrRoCJm4dEITVtNV8iRpCRQu2GZUkEC+dt2ukWKTzSVtzILCPqJy73Qf1SEhN76o
QffIjNwqTrHGe8GpYGpRHS9kFDxnO26ebWgx6di7Vca/UHZmEB9MtFOI4+5rWxR6UCCio23bT0so
ewN3XTWVLFT4F+csdP6OprTCY3g+3P1SuiclgwqoNAGy8u9jvSYjWjQI4yQHN8msDseLuD28sk1y
EvYLps91si21pdMITbQJLLLi1vsbQQu0Rsqyi+90ToYbM2452dce7DZK9tEaSx0TmRZrMpQmFNID
vp4PYUUcCXM2TeIGn345u9xUnBxD6J6UGIMU4JFySUoAbrh4EfYvDcb5wRUiC3xOSfehUY8LAivA
Dy66LkDeIKQDgqAzTS2FUYpGzk+/iuq53L7mVAn1sL2CpgYdSpKKGWTbWRBeGxpBrwfwBI0mFyw2
Gycq4mHL532MvyQMEwayfggFheM7wHXhJLyrnK0IEhmiFL65AnKEE0jp1MVPINlJwCe0sQvE3z5M
FEIf72IW2WL5W/0E5PLj0mS3INgpcmB3rsHF0M2Iltz/kLJtFME2UkGIygwtQv0rtcWti1ZyDV8Z
AIiN6GFh1XHzcuCocpSMe8yZDVpB2oBJLMZSA5u9sxJ0gaa47YynxuJjU8om/wgNZJOvBUQd91Pj
xz48Mul+072U0tgt3o/vxR1uTwpU+A2qIEPORuvgJ6zqhbqrFKFkvyVLbw2BTo3cXnPRQX/1mcoC
TmcLjyEgCcZ7xbqIPyfN0sT1eQjZReD4xcLXlEKPuQc7TNjgNAhXZs6akUmi+HdobMUyJCh/667G
N+ikYnhoYQshvua+wYOZMkHDxOXGEvtK5QNEVwQc8rN5e1waQXgLy8b/w/PiqwqQrCkhsrNaffRv
Zr3YbwlRkZUNCr0ldlyhDs5lB+EQQxYhwsaMa5bwrTECJypS1dzmJZDPZImsAadTHROogG71t9R8
BwlPecHBYcUUDvJxt1W03GzSIoPuYTgUM/krS9TDuK5Ft/8+nOrkYrQIvfdmYLwBm0K6V4jcGueV
gRZVSojNrGJtVFgntI4y4F1saue6GmXnTlbdUAKbgI1aEVfw2kCUAmtIqU8/ZHp2rbGadpCZkNV9
seScLALq8Kdi0TvI13tjhA8RmUTAbfhaOL14q+rixqulR9rXnYr0SeOZDx6NMjw3dOGzCBatRoMV
exwtHJuZAtmVc1k0mtcOXFt0mC8wNl6LEf/s4FwJldO7OY9Wo0A+ocJuJqHUow6GbHMDn2iYvp9v
d0aBJLdZOd9LWVlNcz13HSdup2RIiMMkb8YgewQElj1MJbkHhMqbgO62gaMYotJ6sb31YZVzloP9
OjlUYcwlmmLNjOO+IMijUaYC9DZvNLz6I2/Pc+Dvf+ImOnYPYfQ8yjCDQa5E34BErS8fH8toVCuK
llqy1PmCue/9ujFhPUXv2Ywv4Uo6vV4SwCViPeZ7BK9JVz5BZgjwLD2901mRHdhDacrk1CVBvJEU
FfsjXqvJ28cfWCuChNb3zYqSXmgyMygAY0h5eXVKe9sE+xcg7tvAwq8eL6+J4+QEuh+KSLy93N8h
r2K1He5qEUVSs+RBevY2JVPt/nMNRJev8yb2kOCla5s2EWO3nrScfv2ystrUvl+VfeopSVysSX+k
/yGdoRUTkwDoZCMZ5yP+gG2W7TEERNrL/RCYG9g+QdYQcHNhpnkbovumO9JM/h/H0MHEcRNz3Lsb
ghYV6OpyYGB9FsGiVKoZ/RPLPsXgLoSoy5GkzxQZxJ/KpG1Iqo8Zem+bVV9b51hv4mjNQcf5esg6
xteBsKcMspEEFfQ50FO28GZyODyoSNnAofXtxi6PLM4VNTd3ZGNGWGLPhiwjrPLaiMGMOCLBqvjQ
VifBkgGkcKiNfTJRzkyvZq3hC3DnkRgumv6iRNLUDTgDQX3o9Skh3Ymevd0cAzxAKpG9SLTN8CPz
nDpZP5m7S3xVauK/t9FZC7m/IncG8ZLpF+iT71V8lUWRiFxYetjKWoQrVxxp35hq+qWFpdlwSK7K
/eBygHJbD5NxcxEDG6tFY/NaFZ5CLlCWClToNZ3RsL3yRE+5AEADklBv8oBO9jLpqxgu3jjm4tB6
Vfa5b/5tk270Jvjf/zZK1dTVFV/xPhuGLR5OEW/CRBU19nDsduD1sZKlqpUzRnawSzA2+fUvQzSk
MljfWjSdKxJ81pMGcFV3NBvRNnkNwI5lc1mwdAhMysNWIppkYFTABXozVFNqL6HOR45HBGfXJMw/
GrQR4hkR1NA8/YNCKdokggcgYfrkwglmOoy8Hj9incCgo0BfcpS6WvlcCJkQTK9TvPfyVFwzA7Tk
MvnKq0F46VYpL2TpI/w7FkNoGVL0/yn3ESToC/6tUnK/uUBGNkVI2x+UezFOS42n03KgJFcPyfgQ
W56UVGOkha/sea4+ki7sn85/hDkNfV1JSukKrGnr1fiGAQfJwkQaNplE5mxPVdb46+nTXQaZhuZb
7fmHImDTbsbK11AtmWnecVc6dZ6jSXOm+3/2EYSTic2nHo/e3owPqUKobDcWt3SrQd0obJ+3ACxG
B+QlGJX7yJRPDFKAsMECDWTXh1ezKs56QTaH7q2ziBDgLtfJz1zu4u9PEx/XlIkFGGloW8eXqOih
z61iHwnBP5EnlLVQpMewxz90+lCpzgNx5oKBiPEh+U3J966FbgVaM/7aMrn81H7wLKzS0qbL4Wc6
eMJZU7gXpK5waJlCAJi7g3/oi0GL3xgP2/zZw/QGv6ZjhvRheFqvGrsYRXljrXDw86VXXOUmGYEm
oalwyAm9hLFgKUta1C9uVFQOTeYKDQLMHvaSerEUtVo+nxqqU+P4Fs4/I8Wcwn4RweIpBA2FuGbQ
fu4fzmhLlFvVXk9I+qsoB2lkyx4sXxAK358WSj7yVoK2J7pF2C8cu3v/Bz96KCOUwBe++2mCnDaO
KokEKThNFjAV3vD0Yu3P9gbX2HsoLFaez8Na8D8f/TnXSbLIWz3q87lcUHNy5pr7RGAYMbwkbvID
gkWeAwLS2dqyWeA/A703mlMPmRDeI7WdSWEX2dfIn3M0u9DntN90UvgVX9pgGJ4FphqlpYMEiIP7
pWXjTiI3PnjvORTusnaNGh6A9cMccFGA8aFHpcLIO6Ysje0NJ4SppYEwnWjoTWS6OqxM7ZLIfZzm
bVK7/TcLVNsJGkrAvD70rMj3dd70ZikD9LOA2Q9g9NcohS+Y78NwoFN9PnZ5u6cgyJwZ0O1wcB/G
li48CDCiISCEYc9HKNGJxHgSJguwUDODX0KKNzO0G/Q9Exc/CWFzm+lcE9Ivxt0Ptj/WmfVzsSN3
+DtOhWuyS7/7uufyLq7EubR7EDKYibp+45xPv4y9ifYk5uH4AthcadtwfFzoXv46/E8gamMFH3VA
YMJWhJpSMN+HkxdTGM9K8/0uxBGApljIa2a8QRYS6DAmlCSh8YANe/U+dBjy2lXgW0rnstnFmZnV
hgOdQR33/CR8AbfX0p3BFNUUBkPupqXY9/jTLQNEN6DQ57MkUBPHYZfbCECfrMulRqq4ghPtEvsq
kESGl0lUXgfWWsp/nA4n1GJ5eWR/jMQrArGXc91pwWvEGz8YCbXbUZiB7fGSzrSmxT0AKTEaupZI
qraR6czymJ8cxbu1uentZX3SjSsXi9MSa1xHlLqUc9mCUzZe+tH/YfZM6IsPWPV8i1vnj/Mh3Fgx
wes2pXn/P5Dt7ElTNii511Pe4vblEApbvjE49zYh38Uk9qwhoryohAk5t4Vk+9WXsZgwAOYX1gt5
E8cEx0pPKyCG0Kb8QgC9/Sn4im29P2TeXRkVwOV4ZZVYWpGrZI4ZWQbkX+6LuJeqi/fH5uBxT42p
sAwIOu7c1C7KY9lpCWiV6EUZNtp+BvwzxnZy5Exy46Zu4sWwoQbLnuVHenYrHUxu2hzIDqS2+64M
HEhmGhTJvwB1Ik4o5UsHSZTkslDbsunz4WhIV78+aOg4H6tS8tne5Mtyjwb17Q1HFxpk6Z3kNzwO
eoQ5i+wcgCiBi8F0XKPW/tdgwz+k99l77bxnr5hRo+ae1/rZ9N1fKGPK+ocehgvOBfXT2ekf1I4O
oW6J/ehbVSFINxj9c5Jypw42AU72ZuA/yh1P0yNhtbwJMU2ZSLRIsxlMRS/HSXsQR1+n+TQOOUtH
rvgzDzMeqXqRyDGsanBKkiPEjVCA815EQXDmzF7m6nQKAdAZrBKqu1gsvMhz8rkJon2SpMAeVH+I
4qG5KNqhAq684GIKg/4K7Ar4wQzRPGiOZUOTJutZUNKwjh7gcOBdUTfDVN+voERuDNS6c6q1NI3l
r6zvqwwkWJBNHRd1FLDZ5MoJU/r/Fvzurfmt/OTZwSETvpwY36XMM7FUQVOl1kPZdnfMG3CQ2z1h
Sn0V2qO607V2ziUxtes4kMGmw74aDvcMCQkgCJF9DDXtLr9K+YMt/wW8GtXpK6ISHXpMT2NLHmRD
XsPiY7nFn5ZYh2aYJf4PXV1yZUNQLyKWTRP+tf4WycYDnYSatWSDw7oxnY+vnPC9JAXeRpHrDpsP
zZwypjC+dAFFTTOloaC6sBzXoS2NOqLH9G12PACd7+Es6x+NI5jQ/I9VLzeY5uSUR3lsF6/wOci6
hO+dzcKlvqN0zFpUjgXmxA5/piGQUVuu84jk/JDIgU559jjvG/SAfmfNP8sl1511koZIg+33Yh1r
GVgsURZcXggZRHZIK3oLWvBRhi2KeOZ/52Qoy0VOJ6U9tmKZsT9f8Ty/uyKS7YMtFuXbzUfUTrAH
RG3rOsmZytW6k6+jryr2T1jPK5XumpNY4cB8otK2xdtoJZ9/CdqD8y7tUJo1YUHkXrBYmiJqyVTQ
PGWLXq9y8t3nhxRnTee6V7gwbsS7dsJ/X0nDc6u6j+R0zI0dLTMBJim4hbsu3AAROzK2LzlVlg03
G7CRAs750L0D0YjXxp9aBUiW3McYyFlfszpryWlX+YRuY+yg8Ton26o3msURv0jhIsOLqbperPph
7HhiGFCQCJ+3WTt+1miQwvpjw6t2t/lu6+VudniLPr1L8hznmwaTM2TNbuYZGw76qLi4Kc5WBFSC
c81nCMwdalNM3B3dhF2M2GBy4HTSuWD3BwYpDEC1XeQuNyDOgbA+n44ny2ePB3Q0HgKSrE3Guml8
EWhvhWi4vhnYeKjMQO0i4ADsQy055dTKQ2ZmELSA2D84FOqS8kQ3KSqC/uqHCrSqHiEenSeHy+xQ
q6WENLFpd02/QkPnKkrTmNK8dD9G3XXo7Vx4kzBr7vtiuuI8cjo/SuTpEjeMB5k3upOsYX5wegKs
l6RD1PF+TJ4cffR0+Ol+L4oQY5nt3dxhQ/L9+g70ChOtFr23X+lkMgpygYzxx029B3xvXuahW4I2
FojFaFeLiT5m/kpKW920v0fL1yxc/QRfQXu4OO2ZqxjhqNJNgWZeKRYhFuFslBeXhxOE5EQxo5ha
zpmJUVq+H4GT9n07OhiyIBxAExy46knKCydNHxZMKSwJ02WdoCi79H2+YsY2gVLAp2UK2Bnyjs4D
74cUun5qg4QT2zljd7PwCSNbGULqA9VJWgzbZfVAKN4dybaFQib+Y0eIHUMv1mu08FtXZYBl0whC
/nh8Q9DF4M8rIA+K5jKlJvbNjqXmnBcrsBOgx3tX+pex754q/zfMPbz90eIPJOK5JkUq3TZGMWT9
k/HPPtmzcVAxyXICbnc9rPIdZGCDR2CPW+rd/8vKGu7preSgmKqFOMaoVVFssuyBawictGDvU5aH
Sm7Jds1F2AG4F4SvIi7fmulijpiEov6gMeCniKTGLDnvhG9OQGHw2uvORvDaOi2xW66l2OjoJTS0
sUQRyZRt0CKCj0iLgx3BR/4nzy2rWjlHyH3CPCU3hbD6D1CgVrE8FhpfFbCwR1vcFusGCwXxj1pK
FQlz3JXjb4HYNBh3FvyZb4fZ5UnXG09cyT2fsL1GEf5SxlL9LFpZr8NqjU9cHQ/9EypeJVCMBMVw
k0ene16P5q0kKwp6wT/TKILFHS37fegInqlqoHPLCrVlxOnypaD8eyoDN0MfVXlsJhryCpol0CAY
0s0NnIkNnPezUe0CqGYxCajFanHM2riHDsyFupifhAoMf7wFEkzJMaC354W+F6geagxu3L9jsVDM
UCLzA1q74DwiLh1RCot4ZRs7TEQb8q5AWXyErrzL5fhFA2N5bhmDcu43h/aU8SY/5CnrIoTFKbf6
JGitXYnpOmDTJZj/37cQKLgpOoTUsHvoHwqxEZgjYFipJg8Y1RIN45sEoak42Umnfd1WLPrEr6Cj
Xew2r75Z2Xn03lpsEXEsZ/ZbrjMs7ljT+8MaiWLRwaGHhoUGrKinDrLU0hBLgUTaKD8f26yPY7F1
Ildo8nGCtsm/qD5pJomL2FwjWnLogbHC6fTSO25+ZnZYIlxWmzu2U+J9UpRUPuU0WAf4rvizo3Fl
lnYkYd8yZp52ZNmkPWpzOYR3qLrb5vzVAGzNDLASZt7wGPfzJ0sweHME7hYXYVmzpBuCIj+HPeUQ
JEuQu1b7JscCYl6dFz2oMgbYyZ/zKAfYeIKFfPSK5kkhGxE+TJJjXgKeePAOF226lVNloId///oS
qD1JWHeuoj7QSFz4fhx9pxiZYZ9ZXFmxlrcRedle/BogvrUQvH4HVnKsXH8mxOsRN9zHr9ZSail4
5bWeOr0KPadwzmQlqQeY2WC8+oSffEdbXsXSQyGerABKherc4f5djloNuS/oiIz4El+K+fGx//aR
lqWro404laj4TwlJzOHqEPrnhBq11yEcjUrjp0ZfCoG4xFXeajPIlncor6ZVynBtSHe7riguAxqK
XcYS6Xa0x9x0cB2fspYbsJD/cfykKSm04wQSLe2CSkR1N0KUtcte1/EN8RK2TCONfw9Yc3e386f7
i2RzVd5A8y0LteiG5HJvl9NVE3QDiVH1PIDOuGNa/zdRczlNq8MZxUXyqR5r+5CIPa2mqiDh6v4n
hrc4OeIjwt862HZYYRnEGbgFXMJoF0zM60Q9Fh5P+pyiJgt1WMKXUFtd4kOO4eehwztkOAyWLYol
SKyFI0hlkQxUl8B4vwMj2M45FNQbgxv1XncM+15aop9bCiNgdmcg87cgrXWSxKr4fdZY9bIfW1bq
+foxzuGFQ/FyiAd/2tqyaAw0nxB6sbaa7C2imChiRazEFjT+z6clLa4schtElK0QOI2rpW0lXUH9
ArmaLATFzqN01KPaFH4p9/CQ/EhZCNBtkFMULcJc2SEAhPjTAGbiHCYpp2xnWQ9K8YvZESI50q0o
k5mUwS50LHPsOiVXillALY7ybyE7gMmGOYgmNmOI9zhvNLmt6QCrVWrEidmrOj8rROBgTyJZ/8p3
EAP4FLXfELqor4ZS1GlYtvOPM9cqxSfbhoUqJ1ioizHRNKkhetzisXDlylQawgj5RMazOlqsLhEV
FgWJH0m30gA4ORRD1m5nHs1rQk72nLjmnynYmB7Kh1kI50zEjzjLr3oNUOWlNz4S8+RiYmu5Z/jc
25tx8hlJbj4+PC6vAz/cPl5aMFYb8MqwcU4dkEYRO2DFNWaCCoouLkCqM3PAiybvo2GY3NwYS3jF
U8Fj1PtJeLhv0UrxnVpBACppVjD5a8hPX+XTWGSt3hM5XP9lbDIEiJ7wq7azpoBd28mLGw4BOKIJ
+tYjAQpLmo/2lNEY5XjJIycsCs9D94f0SvdVbxbNCkyV2ni5iiQjpU7m8nMy/mt6iKlHIBWpn9NG
KeAvG5FiEBy3QhS6vWTjJG535pbTChUbyUIkEkC2GxhfHMbrRQ4DrCV4mHLA8PlaDz5iABjn6RMY
4pj1ouLTwGuYK575Yj/R36L126fHnj1tzUylGFS2/xpHHY4Yfx5v7wnRaM+GBJM80ZeJE7sfVcwC
8QeTPixF0NAlRiED5A5aPzoPrY2402kVgM4214704CK09k4zzIy5jjWXeNjffcWEVtnezx+YrxDS
11hajbgbfbeB9LFslEMdMWU32JWxspLrkY0oVb2HZZft1N0N7MH17YYS92W/USJBFTt8R3O4m4/G
mtISNKraECA9kTQKwzE5qoMa00YVSNUGgZowHMbFVVb9AbDtQ9tbaV5NwLyOEmBrurCUS6KsVbG/
9NZvA6GtNIrFa2D6dUIFqPwhK/EU0PfJNYVXKZ3qRiLSne7whokf0bk5eA089AYUA2pbbI189yNQ
V4gw89NsLM7OWtk62XCQ8QaRpnJnSUMkYZjLnvsXLxM9ODWxnkqAe5bvSBZQxXP6l8xfwn1HtJI8
RFgdL3jH4ZaWaEYHfdSfKM7ipeux3Xd90YyPlx4ww1J3Nbym3FWycWBhRWkeCQS9R8cnOfFe7+l+
9zoFV9itnhDCoq3YDhU7L9KcyRy2UCZdUQtaqip9GeJ3c1iv0aU5pDbyFN07kh2y5bun/GccS9tj
emBsVIauFWDPnpVn8molzXJ1JbmOKxICOs6NwZC7+AZxaZom1haKBFrYOzq9HCKu8vIpUh9il0q6
Pw4rEU5dL83hDXHAe/vV+x2nKPuJvddFWYzxVolR1qaUY9RtGyN4lSZwx150I1+oWfDH6/mC4f0n
MOrBzIte2OROhuL3HnqGntPROepCXbZBxh3S477V8VZSGR1pVy4v03ofN8gJnXl8/SGjjCKnDIhy
ZJieCvI1C43ytlmtEgzaY1pMr6ArzVqdzhzZiI3hKVLS5TgXM9WjDEwaJ6riiLqiolpMWhPQFHiu
bavAoOt21cTJ2wYcsTll+rhwgr2hxMmznD0RLuz1AsjGEeMuUc4U8lpeF5HrKSP+SI7wy6ndqFnJ
4beEmD+N8qJeDx6lTU7uhdg1DFTHDqFdiA7xTuq2d9KWzfBRDU8OiBOpgy0/vH6uiQjQtfTlcbMa
3p9lYZNI01DPgjPG+Dp+Ohe52O4N6QtJa+gy2ChfWYEuNMh8zZ3k7c/F8Qtq2r64veiYPDz5Zwpr
ItDbvNH9VGyxfZ0M0znL9WpoE+YvEkOohrXo61b2eGVfXbgBY+H0WzkbEvxkCDhrllfgoOdeDrOD
WhKRXZVfeuNQqVHVKQomu1Ef22Zlb/Y1/m/H+3eVgEU6rRxStnqdSDuWvLtGLsjqWzXyuwBwyg1R
XtX6HL0Ctc/2zPZ8QcZWpAk4W7ky9T/juk16bc1C1S0Mbm20DUC3eXn0+HDlYiwH7hcYtHgjeXLM
DWNyjsyox2SD6vf6FJgnswZxMoWXOL+Pd1ATsMY/333IASIi7iF3b/USxlrUlxV+OE1Pk5xLNzyU
utz0UBvBdGqylCQiu0uHgimR3WFisqSmbftDLBy+DnAR7MPGfnWmfpmioVlXnH8dN3NMGy21ysx8
JCxOevtAVVh6qeFKwsAUxgBvamQ1msGfyCQvq18wMFvKzl1JNP902msfckh6Nwk2Un4uIgw7rINv
Vr4iwYKddPyrA5SPBLHAA18jy3Ujn6OQTLBP30FgQCR0en9cB5rviieo+yntca9lbVeTQRh3kJuG
YSTlYv6JsEMYYn8jJg98xYZEcdwi+vrEz+gI7GJUtn7k4sLfHstL6oN03WgMEuaKKFZtLpPS1Rbr
/lJyUZ0lLpCTt/3cJ/K/x3mHL65SoBjuxlw7iZPSccpIIB4yBA3jGNy6qoNeZc0tTiW/PG4cdPpw
hEkX4A/oWZCmdx7mGFrf9plzg4ae+W68Kk7pQ3TtI793uguYTNkceQtHZ0YqRcpqx9lSl9bCsItM
fUo3bTDAeZ2tQKpvPmPBiLwsQxrAYvKXLfeuuc9jKqqwMJwzI+FJBlQAd97Z9uHsb/xWo45+7/z1
e0PGjDaqE6C63Fokg+rKvPiiSqn/qDPtluuTyK84QUDNS3S/CCR6S64QGO44ae8OMoaRMnqE0jol
WUq+PIB+0H2TCq36jP53Wj3kEL0KOEYeEEFgCOjO+HNMMReBslUu0wEic7sSbH1fEDvw6L8nXtYe
mLHMQ2AJIaoJXgBgtbPd8+vGIOvyNvcImyFjExfrpmIb+5i7pywTMgckrbUZFEt+pSI/TrMJozkU
i8rI6boihGBfDmu+ow58Vp6cKECwOXNmMEqqTYQ/gOmA0J0QsR2XQWKoMD/hBFn0AIlv1d6Eucty
WT3p8X5a/MLgHjpFsLM85AG8KtwHgm/VDcFxrMHBkFtHLw+PPCU7kEAJZFerVRaoEfb0ApBcfvw2
UCTEVQUB75zHcM/IDJUxaBFdh6oK8SIU0lxJ/ODNeaYQWEum+khihTLID52YDJWshupv76+pz9d3
8NNs74C0wlxufV4mn/2GKmjUI0CHu+gRU2bjgxrzWU6ppuMLO2kWorlU2SW3UXYad3x0epfzN0B4
wx5sZFpizCDqUfirjMo0DpqW0zYqjUUeLm6BNjWqvsvqHY2ixXFUS4HlIMf1sYX5LacHh9wo2w8H
tJirRAPqli09a8OsuQmpOUmFIcQNUGCOcVIadUZ9m+0XQ5fhjdd6G83Zh7BYK5qUSFkIigGT0pEz
xO/RQjpKY79JQladT1R1zFZM/xfyT8ozuwsJgz5IbqMEgA4z23iOL8SGCNC5irJoRYd4KfvciwIG
zw6vaIN71gnRqOJQAEWrlKInOBQA+jkn1O1/ivbG0OvqqhBWrqUZbaekF3M1s05s7DFBlMW06KFr
NQU7JzvI5h4G0zk7uZgPFHT2YaV/EJaWPPLM7oK8cKhADjZqWkc5c6Av143wq0I2Nke5hUOTBbQr
uIuva65dINpJ6T8zUAXczqI7F+OzQqQyj9E5Qu+upW6ipW0LHEraIaz6Z+ThKnYX6CGDcsDcjwoU
7CVBUlUw7K0a0CrQgYanSoACBSSddnQltFwvucHQeK5Jr9pCzTn3H0hPn1WTwetbvhxbCBhFHiQT
y7rujD7LkfbG6Q+YZ+OY0sqoLvfGlsnrDyv19P2TX9NU6257jv+Hv4lSl/y69Fo3VjXCBKpFRYoo
tn6LqtM3PQlLHloapQgSUFndeKaEbN1YNnyqQP7FVT8kIcbHEo5Ko5ELTPjdGDHHT92mkitNmbFk
cAxZTKymrcV73t9u/9cxsafIi/GWPAiCtSizSjByMzGkdNIjIqbKqRU+hL2wFfHoT7+X7z3puN9y
ZaEcedHCeeYd1LWsVWWryIZvhQQ2S28yAZfOV6vDi2etVtsLujMZzrEWEJy7PAUvvFCI7JUlNHjv
DvgOcJubA+iZREcGKsSWYR5EM5D5Q9+xQVAs8zq7vBDt1KD2uIgjMKgzWIrNe2WBXvMrNh0XNsUi
Z8HDwoXdsCmWsrjNgaGDOCz4o0/kOPtbvFooGcvIrR02w7eOLPz9WZvgZr2O6lfMZhTDDZ0x7dFe
/J6eAtd8aFaJHfZLGRUfnJkuuGm6VRVArrLvyICg44AQ4f1oOFPHGSexjYDwwg8AFROj94Ua+t7/
b5m0V2t96sV26bTZQvRV7Xaei7PAc6Wc6CEcwXU0vI4Q6lXLkA7KtcW3bR1+blA64vmPwX1cVhry
RON8ClB25D2NMOymgqsM59GTLmTcM+HX2N0U3UPLgJ8FUUn/UEAR8IKa6Xy9yRVf33F14TOBUj6S
6S2DV5LMczD2SiTak4s6I01jLXHq7VFKgB+s+2advo9Q0tSruSh4njYsS2pdJu3hhFkSFHuKfy3Y
RA9Z5XIZM4ul+C/ErNBKxb8qmvvF6coMj0on+TZtNcdcR+DgQIHRowxkNSK/gCwEC3YxJKBUwTUW
w5lKBe5W/ay3TtJCLKk/S0EfiLSYAEyRztBf+0aGh7NsUyZpeXzA9OjnY4Nvgql/mDfCqzeNaexD
hyO9Ns9/UvYBV/LfjHZhn3DQUH0F2G7lFfUs0z2jjtv9r4q+XnGwPOs/WPEGtz/eAqExJ2dXxCph
0sGM6vkP9hwHoa+KeSPipKN2Iua4T/jfLVq5PuwzL44qbHLN/rV9hxKRRoI6oDrymzFYQrjlrj0c
SqhEmhsi3FFFqPSlKt/oAZHt5C5irwwasQzns03zHOwUUHvker+O/5Vlik5pKPfZN+Xm9Ej3xU7A
Zz+d2CqOpSlzA8E9trQHLLTeUW2znYIK85xA/EXwRxKCqckt0Bq0XfwlQpAuSJu37Lc4jUsQFt3g
DiLzJy+oVjEKlzhwlAoQmxj3Tq73m2GTMM9IL9wwWevMYLPaEpDYq25IvU+LEZiZt4lqanRJha9W
/jsBEc19rM5HmslRj66vgOatifoRqnnbSilsztA5at4YX4yndyaZvm6MXS7osnEqpHOsCHN5a5IV
XXN6/iD0AiKgdsS5balESsQkv0eYSOF6cQzeKRRDiKUHKeHTGXwZgUTBMw9rfdnu4mthv/qKMs+E
NGRAknOm2d1Vqpw9QDtNDFEzrnQmFNxFjoY8JAmWSL4QxA3nqWIm3KOd4QaHO+3WMx5uiZ/GGO5D
tbvXNlLeH8gC4urs5X2Huz0UcQ08gS9vdU6oqzz88xh6MF+Xcg0kkYYy+E/IM0+IxC/RUPFD88Fs
Ad+JWo58uKIoR1aL4CCyj8a/VeSruCjhdzcKSEeZDUJcObUlg0txGL/gy45J1qxxgw9uPAC/7fwg
ullps+07D5C+JmagGhLIY8nAoe9hVDcXWtn/PONw2wvWkF9990Ez4aAsPnKlmHQ4J+3oQPtM7LjQ
+x16bw4WSaEIIJdPrb6Lb/aFZhXFDrxWPqOzWK2UtT6DGJrAMgLru/bjUw1I48ZTMvtp2NsdPqeu
C+syE1W7K0vssBgnDf832umXGBvb5z0SXdoDuQFDAurKI/4eF9lxPC9XUfu07dzeiaNqqzyPwgrG
djhhmmHw1D9XYNG6MwYlCIXvgoPWfmAgl4vQHxHjn9eZaE+8fKJfH1doxzYyX7m/TlMsUSTzESBV
NgJr53W6iVtFQT2SJiAEiTtW5b8GixWtG4ChV0s91HLk8pai23aUxsFqE7iDKDOTcGN/ZnM+Iv2d
Xpn/nlyde2QKhV7wOr8EeT8jgCPaSkbzybFtz3yU/Igq3Ae33SGWDuod+Mop0oGYrzTnJnT7OzlU
gJKYdP+Bi0Vk8psStifI/LIMmZHc2A9mqV4V7rbs8CIUwQ1XeKVlxn9obZzh6fvQWP6mA5l7XXJu
Naad2t6TGMFzDfw6C6wodZ6nE8nBTmR0L1ELf6eUtNNBO9yZnBdUI0qpH0CLFjJ1zppuhqs/A85y
VtGxWnhVHr7AHTtov2ggRkAQATJQPriOq1oeNzlwINKpVtxAF87c3bQ7xaap+pXwAicN08OsTZjb
Z7N3cHG4V1y7g0nQBLLe9fP6AZY5qPMe2xuORcpFfVwOfpGt8V99uZ4Ol+HJ32YxKO58eAyRXKnq
7AcbNsq1b6258Q2LOUti+AI2H+7YpeJBek4IfFFJ9NW2kbvnJGN9wVGDXjXSPx424U3Lat8En3ba
4qDj5vMdn7P714XJUGJgpvisMP4yXgrwecFgkEz/It3kNlNBb1cUIqm6Xq4LGwCh9b5iphCFpqD+
SPbS+H1zcrZH9XKc0eICdx5D/rT5VTIE+GvZdsRcn3NDVXprexeg1iYPSE+87dzIs5nr7/N6ru9o
mkCyG6ZFJoIPmCCsx2E6GjWXNQFQN4Tp8fpnGldkiA2rwbdmDtC+3VVXnk0qAtsMjOjqrzemNedy
YM/SIlL/PK4j377Ucq1usNd33zJO2tbrcEdSDrkJIIETjs9+wcjeBJ+6fc3QnC2IlxevS7agdw+g
nQjBtPbVzvLpIdPsxZy2lWhZAHH3PZo21fx2qd/TSYkhZflqHVeS6cRziwdcu0XM5pG/sm0d8wyP
AnasT7LliKGn23rTTPGr9KZzz4JNJugyDW4YGjHUulxz6Y/8KHPRl/CoAaxPSo6dw+H/MKGnGP6D
jcAXRR1X0mLcimaXjU7N/p3dfnsdK6KA/ep77oH7OhUzAt26tg33Ha9ms1/NEdbzJpdKWy0fTkhV
2TFHseCIUXYBE1LGvuj8TO34MratcQ/qm3hTM/G3/LEwXbClHBFCrkSV4Qcu+bjjWkvYDTOUEcQY
V9TY0X/mt9XSw9QeszisJtWnE33MilZUd1xsl0AyqgwqBC8iUsPlcVVwYCCWviRZdPsX1UqRycmU
NREB8k5rOinEEkp6R1olvbuB1P2n4Om6NiRR1u5QY69TtOQR9wbqlZtgZ5i8TuWSnYt06PS1liac
d7hNwYf+/1hM5D0TcFFjN/97vHUzbWXDWf8pf68LeGTDJo3Kir6ySlPHRQV2+n2oK6zuA9rRhg8y
p89phaMX4peWfjFu56n1CNHnUeCSD2RVNmRcgzp2UxL25LrxvWN6+PG/5ccCiXVD5qJJIEhoyOdd
lrAv6St8FuAuTRG/ly0KZEXhJU4lYsXZmETvE16K1QTMt+Is464OVEAw/BO4A6q8kDjOJheQnJhk
neahacsnH7ZA7+dRQWfTKAoleZ6YjyupgiCy87mLImD6jH9RDH66r976VynuY0N7UY4Yp35Y9Ffg
1uUBENm9YIxTQqMxeFiGRreyDhbTf/J56r31lpmqY5RXMb+Rs5jlW+VXJ2nT9ZWYtLRghpio7Err
Fu2diWYL7hB+8bo51a4jRYMdNaLoBZ3veMAuw8c47cPKZ90OVi4Bgf6QgnRxvz9B/HPwDmRMzKA/
qA4C49h2fh7xhDXpp3hVbPGp7+w1Uxa/PZEsfzSHBYw1pxpV/DiIgJAyihXbRaAK+1HUvvJku1/e
eyIsLU9ZHxMh8YmCpx2s7bJCmaHCxZro9epK3X8qXQyUaWlpuQulVHUWJzN/q3mf3esQsOcQEP7c
O6ZzQCC64zVoX3U662+Qp49/aSElHOTolzUEUU+9P31Aqc6IvLpSB8CmrLIz9sQhr873HvXmLQaK
tzvkl4xnJjkE0t7aQw75sTpW4EIpGwa8dd1MmuefMtsLSVTNWPfijKCDMtYW4gy+IEkhaKeVLUcw
pYtGltQMRROfyIgDzjYQlMUIaWXXmxX51XoozdbmkMtiqqGzW0sVtv9Wj/Kuwt5VtKWhW5IvD7Qy
nDfTzueHn/kVnyR1PJ3QO4Zv0It/L4YYTWXCZBEFPOsu6jbkbTPTJsTDCw+nCTZmSOlKqUSO7hO2
ov4JGr+jb+F2Gsp6n5ABuU+lLDJQhKmq+ZWa+wbTCV51PO4R0R6EDvglqfjXGeif0nsZLpzKa0wS
2eKvBtssN1+DOKBV9ZdvMJyWxEWlkezK42BY+1gJnEK7HPhOjHUMpRe8RKqE+Vat3eZvZW7zbh1s
AWPb45cMmOWl1QZtvCi7I4AcImUlY3kRyluKTASVvQ4tXu8a531aLBxL047yL/RhhOBZhzFtfSvm
1AriQI7KsfMI+e3WLmx6YzQWD9E3dy9KkrRt1UGcYIXUBWQoYH8qeYkFZlKOGoomxoA5lzdYiNCp
0OnsXBdQ+6h6hUMfrRu6UJDx4rdlIQOHR3cgiyMIg3JamcfPb8KLjyLwcNYW7c4oZPqJaUlUQ4xV
fQ8wbPv9HbPcaEFslfitnWf2ZbiQaGTF95wHKfVxnfR/diDQR3ENPh9yOV5l3imeW1PfN45u7Vni
fiP1Z9kXU4U11Iqoh6wfhQoIo17/5SMP/P+bJoNIPyDEN8FU553MAwpBGibrBVCSqNiRSvSmQILf
gsn+y0UoXYjyGJ42UXW4Z2gB5I06Rp09zLv1G9T60Kgj3NrWvyXHPIMePbpEnYnFLYENGUERsPQc
S15/9XpsWB9NQbScaeIuivaLBIb44GlYTaCrjgYqqxP2nBLMGLiOMoPraDvkaXd3vZHZBe3izIXu
2QOHoepNI4KKeroQ4enfqMWhnNGp2UTmU6YSI7t206AboaBMpE/DqCGubldl84soYc/RxLAdiJ4M
fp3G/uTVI5GuzdiGsb40SIE47AMqJmbc1FhAIaepxCz/Nua4hRpllzd+59sgCpnuGxDuLmPW4yYh
mdOhOmH5dIsxsw0KYafSuh3brhNsouAYkYUqV7Aglp8UFxEvvVPhcYKKEK7TK3Dn1Nmrk58rCXXu
T9Wl+C1DCSc/ckNeBWS2OQyOPUFuhaalFTnmuQkztIiO8Ukt5ZJlaanuAdPVM1Nt27QD7KlJbOkx
UZIzAqc6bghB7aMStm6/7yByfQeCxGTqwIma7UHY417CpPKjGRITZljI/w40xe3O/xSoQSLKHYen
gvz5CML8exkO5/h3QTXEXG/oMDrDTfC5NfxWEjqwmBrp+KemxkeJW29BVdQam2cZLfAbycyndfA0
U+IB21weruV06nLRHdalGlChHb9moBjRkrDSY53DJ0zDXK7rEUgCn13bDL9oYnGWYUDDeGITycET
0JeCRRbq7l3KZLhZEe84qKISXHADZHgFeWYsLmekU/q/RrbKZ0v56KtwsQhIsF6p9+GtNIi7mCNh
1pZbskLSt11nAY52yXLWgI9OcBA8yuAmrn8Q2AYvyQGj5SJOpJGEV/3m+uPfmPQW4l5SmIk7H+cx
Rp/6wIWdbweqo3xFf+ZwIoIdl3MSPTjb8ovTaTdpwfFbo49z+EjSUnF6Y77laIRR7gVVbl0SUoil
2vyCWlvf7PExjy4sMsbvmIQ/X2glBBVqiwi7g78Z/ecukl7K4J43s7xFauS4Hpz9OR/GNDMf5LpR
Un4rpPA+Xfhzpx7slbAjpq+N3CXDNZ7usotXCTMCjAbG5yeek03dPJs+Loy2/yGLnHrlbHYZ9rgT
WR1N4zxIHEeMYOsJBNkSQDmOmAH34YBBwcj6Y8Orgd5fskAA0tOOaV0dFpGfmcfN1rw5Aw4W89Yr
H05iIqyKhCAcDXre3PisDS+5qw60SJ2vOkETVV2ulZ0F+OOK2ZGofytVzABgEzaTfg+go2YJxpUZ
4wb6Hdf64W9F3wJFczryASAgx9TYOrKKHtfUnWpiu6NH1Kl6hOOsgo42CAStvK54wATRc0rgtwxM
6OayKyQweib7boNuriVKJwL9aE1nwI4hapVeSUKoHDlSvXEVoQbs1fkgGKjhTAD95ju9hWYPac0L
POYNrz27Km0TtAqK0w0wbrP0waiMlC18l4NMGrSz2p/hrwqIAcC0y3bcILbf3mN3rwmuoM5rF/KB
lMzlyElUGdk/w6wdT/zgS3Z9Lr+CetxOjjhSfeBPKA0FHjYGnJVVeNdCM41Cg6y52j4bIveWQkKd
PX+XcgZCSl8w4SJfDg/Dy4Q+cCFSAKDUo5la61l18aAeJ1a8bHRdMg7dLLCGqMcwxcvvPur7x73m
L4q1f72MqyI/oQ4diI3OmMGGPvha+byEa1jiEWqvNgvh9exF4OuPugA2k1IuhsH8E44SeEvMNUuC
C070EnjIA7rqJenSyZpKuVnf+7Wx5gIsa3K1axIxbyAbFVJ3ZMgrurlqJ1aBeP0XZd8uScH3mGFj
GofGCgLU9OMC6Whsp1RVM53kHH7t9p6VoA/HYwLTErfXYFVZeS03apwtmGA5DxgQfWhji3Az64gg
x6SmKGoeccmaqnppYDN7GTSHvU+xM0bdXwytQ6Tdzsj721U9aQ4NASxFjRkPLVnHe4fgrum0xXn4
navxrFTSbZkIvOYsejNaLQ2IfIci2qvIskv7nrdbsXMJCyM6DJQCmxRxwpEaedbLsuUPTglpY/fn
BpeQIxN/8odJ4TRa0ltYdjjN3ftGK5R6BO67lBqNJXG/2aKgEf4VNYTOfwW7LMPCusuvRPSL+f8b
eIe6iro1cUEkPjywG1Z9iY0ZjOQFhUwSGd6qHNPLmiB0gFdVc1o7GXeoIKkGKrnOaZjuDJtZIebb
6UUyafbbjKDfF14jKtUFoMLfHxslX6+lziRcTeF02VTXtwpXXTc84dCXhCeOwk2/vUCrH6Qg2AIc
E9Nk+vRLuW0m62/Ck5TcKqQUfGHl5AwMTwEFziHbADvxrEphrZQH3F/TDpOG3CyDrjzluHyH9M0s
L7TCdNTsmoTI/5CpLqJ6YwhaGIybu5WHI3nLhaDPdLL1UmWYmAbI3iRbnFVSdOowYWSK1vSO7IDL
PQLFv73nKwt1H9p9lRR0pmNEPs6IgZdnz0GL5lRIKQUc+E71b7zGmXADcWxdW8JNwhnbikzU1zyd
knQi03agCekcZ2TrKm36PV2rhp6yp47DRvsSmdoU6O2+dQ1ephBnX8wbAhLKV6ZJfc6w/ZTIaxA1
8dJyjFnTSw+VLP1jg2zVa3u3GExesnwgWN872T+M8mfrdQtCUFg0Oz9IeVUE/wW5EHBSXocot8dx
gLtZCgtgoW1WYLJckero7BZDS1I6eXkrjlODM4kqHaRLq64EPNUXp9V7qPoJk5Bm0SuI6WIGbz+Z
BSFhscesh9dyb4XDnkPTd6PlSAE5Hw4/9yMg07rGj+saHeBiQNQlDJfhHtP8MrfSsiVkSdwvhDa4
P9gxQjYGgX4Vot3LjP+3OQFvxfcKOazcnLxxK0rZLopqgKx23IkSy+mB/+ymEDiBgllA2tX5FJfV
VSwEF0YM8nyVvLNkQeGjtU/0hubrrNlVm0AnsZ9aTnbqjP+MxndQuSsZqE2x7TQMkxl5bzdSPqKt
B6viebBnCfADBwzGFHguV+TmloxzMiy8gyiHD3ekbFB70dV+G5KaxunNzeunqXyKwsJRtAf2Ug4Q
tKHUKuDLRi+Sv75+YNtnU9aKYPRYrPU6ked+yGOkiWX7cQspVD7Y9FgkZAs3MnT8KAKeMTZy/ajg
/fp+2An+9FAJ3WxQwal2nGLUHA1PD3/udutqG/1ckWpMwpZvZuPz3LRbOBcnkmTI202uD4ALbkSt
s4HJnzkkARqgS2EpjFOT4C6yB56EvCwLxRwFm3N3lctoapE8OCNohPeUCFfBOPFkh1aKwu6nDGcX
DRbzRNTihdfTPwE7aw610vidTiXpDBwvfklQHUhchb0uAUEGG2eNmPF5uzxpaVomO/nyS/6qp9SF
5aydxq82h0bvfoo+7LkqkJ0e4Rrcd40bArLWG8Zc36uaZeK6St25uplfMkLkZFExF7Kv2P4FO4Wn
ysWnJKkkEGAV8n4XK3HAY7wy5Eb6DAOij68bMq9OuETymJJk2Ls2NruBtpLxruitJnfKcqw9rRmV
ts0+hWt4P4Owg/NboRnj9ekOmJiVhAi8uCkrAC5WQOoRrPALgrKrnQFx0YE8ao11lKnWmtclwkkJ
8k6ZfWx7/aL2r4pJCQbuaJg12rI8Ahi6jF8hKNnWjIvuM0AdV6GK+Ttpv4BAo0iHT/0mFu7sbJaF
xF0kSALpRN5IXSdaXG5A44ESSQ5ceZ4ZOabYeh//iYePjSR3dRO/Va7CJOT6qoCCAg6krLgZUu1T
b4O4wqwBxM/serokGAR4n/EgL1xTl0Ly0UuQuNCZJ0RQow9Y81GFsgmEnDW5638OpHlOkjjxoKXI
NrEijqyWc8KO0/NzQeS7xFp9P4wHo01lf3S9tQT/ybTRCodOgGH9chgf+ggVIKBvxBKQu1vp65uu
oW5Z4GDZGfYrUgGmr9HtHRozm7XWliZZbDcwC5Tduq8CkjWm+Q7uHyOnAHor0yN39ohAkb8h/9B+
QukLwy0qsCRsUoyif1S6S9vToNJIxdGrpLZUcU/y3ydO/tcLqZkSEDt+V+27yMRD5NHFMHFda84d
alzBpJk7cwkKG5x6zlYFO+E0XwippkTGnvfGGeIe6nJqLh0t1oPy1skAAR9tYeveyoCTw9q8V/M1
XV12/g1ju+8dSZDLPZjKJXFv5g9SmdE3hxj2RINxLQEU+OYM5dzxFrPFb6YzDIbrdRvx8GnbkuDE
VUACvATnwO5itqraNENPgrurkyHIe2G1MiGPx8A67L7GFYUaJGuykYMSQvHzHY7lbkbWhJUYbKvb
N07jAtkbDIxvtaGNi8WhT6k26+J9zmGFefSFqXv3NbkMh8R9BJOSeZrlO0EiF4+FGJCc6L4dzBbh
4mV1dYIBd/m8lm/o7E4GwKnCBd6lp+WFfGtUe/h83+BTmSACKGXgNl2e86on2ETE8iiMMp9saqSj
eKtjr0YWzTyKqz2e4kRMJeteTkWOZiBJBjuU4wlzUW8Em3bbHuq+fpi/jQRq46PGsWcapieXYDhm
dBN6/bc1mBGRCmuevYzTnEL6xvpCoN/0Mxb2/fxzx7KUN9DqC0nfNmWWojRKeu3zUHlsM3AZ0koR
pRle9Z1KGYCPhuwV3b1PwmOcGmpJlQQm44VvcY2aP6ZEc3pDzTJn9UlItD5of8QhJw6EEIOgKDw1
ug+Vv3onq8KNxwAhqR0ka0TWcg3duXyFvjPv9AR4ZtBDnrytoGg5v+ltDQckjIiJ6mSnWgv/NT1C
+QtIH8VSiUwEDDrtRSdrxMiw5cjcWBNEXIdTAlPsuFVznkkeWR/NuDO3Rsn4HLd84zdZHPLDdPDz
Y7tNSjWgx08TFzkBnYns5CAAKqXCJuiik3pXP/Gunh1aNGcbCQc9oHTlNzptOiMENfD/NDtTiIAN
hXARhRMDOiaNoAZWZ3J/uR2gAz01YwvHA69phCwlpLby3O6tamx7hWQOfMlq6plciRbYzO5/T9Uf
dflls4elPgxmHtT+UNij6IQpfxG4z9li/b6hrL0YIhNvmGmRZtIYvDobNdEyUu+5MM2zqffa24N5
Bzaz6nqm/sr5nQt8lSJaaSyDYuPBvtyDhBUya/uvkHGRbzX/nx9/u2n8BggEbzVZ3m07UTsu7/94
0wzBaT40X3LoML0BvEDxbpPJSbqZyJQvVPx+MXG6hHyN3ANG6RZNc1dznLxsqtU583WF+4F4jlts
nqzKC0EHoaeJpqOso39WtWw68Ui/n7IIFF6ROX5aFWknu8W7Upu1Cdt8opyFeBB54x7zT9q5bjNB
B4GkYjpMZxwfrq6qkq2o7Ulu2wnu4EelfgXzdP7wwga316S2zsnNgHwfIc1U9FyPj4BIhoied4kG
kVJEjptxXEgQ6fCo2QdYz90zvpkEB77iAFU2nLD0JCGO32pN40W9SC6lnklHEBkTUyrlLGZvhPU5
lEbAvQEbwD8o1mn7lW1WrgUiwltEIhqKwHkMWrXz9OSKZrFlGsIGMEx1Olb/0+RHqCiw3Vohn2c7
2NHx6N5yTzV4TOGaPGaavtEOlRDBCE1YzEfwKD7TeJFOYJcbyu2N9Po5Cz61idU5PSQsVuNLX0EY
YQun4XVNGQBAv82P9wP8XbzVExikoh4ur6q6MLrx3NX4gQahzenbOdg29/cZycq/okrJjNJySQcN
s9oRgZzm+UK5/GmameJbls2kwkPT4XQnBQ7eC7n0m4RD+/+t38VIyFSC5QQDTxP5tk56LLWg/gkf
WrLc8FIN4xEBNpzZa6LsiqKxzcWA3ujf2xiwIISj5OzFufVqWpd9x5+0brZhVMDndHrLNnN0zm1s
U0686LUfIl7UhObbs+bikdsMwwlgxRxmrwsDxi2uHaMmkkodda8pAPAQwT4ZMXZ1U08pkw+138fB
iyUMx4T8B14hIbB+5zp7BJpUp5k700DsaASoVaZZf+e1Hg20MCt7uRaqb9peam8kljz2qPbQK2vb
+xJ7KmDQmwAvVYrGMAe/xRq8lClIKWOAPjlyk23NKrdBqbwdexXzx4Pw4DqI+oFkwt01wavTAlgF
tsFmp+uLL0tQIQC8u/HlUgbB0dPpTNym8Q7sQ33/aaJjOAMk6NGLfVAidubIvaZUeohG5S5sNmE7
TQswPnJcRVDZL3ss4tXjrX6zKcNevwrd4YzIgIbxLo3rmkbj18j5QcNZHQ74LUb/P6tWXHxVUQEz
7YFBjGd58s+g2ggyfLhL9FxVLubHtjxnBf7yld2JjNDQx4HwgPVHH3052YNuEjKQWctIDLRvm2W4
kQJ5Uf18FRUtKE4a3PmPk3xBzWjvef8/xsZUFQXHIgpp8KMI96s4kM3sNixjxI4TMjQP2QFFyRa7
N5eJD5qPIE2AeYoHaJGNbpywTNKqq8aVGUTs6uienBidwBXew7QFfMMkxrMXXuhhi0vfLHLkoSDC
T/a5qnNxw7XbN15GzGeIzKTxwPo0lFQpNrwsqluS+w3LIkSVmBe1MPSuVRZUP8rxnqYaFAlSHcya
OWum69zfJQMOabVxtVwxsoPMn0lACr537cIlfw+OWntL3BJXyE3mDp2vr2Gwts6Ah384/RGUgHR+
EGL8gnwsvP4Xaenu/BFonLXI8gUO1Uj7DPHK8Uj4qQpMIS9wscLfwybxTiJ/8FR5FfW4HP1xBmEK
Y/jTzwjeTVFiqSVHur9wN6DbnJ4GIBytRiE1XaQmY3Z1T9Sq96NiWbuEtP9DJLQvWyPAoYbb1mMy
WT6IReDPv+p81gEbYd6LYfFYL6qeal9oKAXkmznUPusnlLssAf0uVkkT8disUbxtlvBI0dGQZ0gQ
OpoUROho/JxR/u7WprC9Uo/hkQTl5iKPlJi5Jr7TogockbNqD0a84V1y9GQsNKjYfNC/FjSRLbcy
wMvzNGgjkvZwbrpSR1kKyhFEkvz7dv2fheBfOtGcjAw2GQoD2XBj1awcPbcbvwlGOh+0KChIRzPG
eeW2WayA7SisJwLXPXa0AZHgncZ0KBUXEBKGfbCM+TlDnyUICDrpMvwdSr/xp4GfGIeZ5I/WLdmq
Wb4r17u+TKUDE2WByyvKSqz1/5cAdZbhQmUn2jsRGcTGZlARqZJoWALdD9OJgtLtXXdQbRNleBJ+
cOP9MfVC8xyT6+1KHZa6w+VE4S9sC/0tG1vUgheWRwqwGrZgzgoUcwfmIKyXiiEDfHsdQ7V6VGi7
rCMB9QLXWhjI6PNaX5Fn1gqy1Y9sZ6Xxqldj8nGZdHzmDLgrVOEso4H57FHZNfo9fFSvY/LTT5Vh
ZvjM9DYVPh3WaJ7a6iMR+rTFHdfoIGDZnCQxe/y/3pSYhUKVb0w31LW5WrcYoVD0h6Qn/+D7SeNI
HyOx4kcrvoY6wrzHIiZGyQQTHOVyGu4mJBWKdXUukqxZd4wbxQ15SxuBPfriYwTqr35Ohg0sjbbv
IphKWQ5REi+q9nKNsGso6gvtMt7ESMkfO0LuikNkz88itr6N9IEemExzVaRINyylj/Nifdy/2aXq
RUw6EYyzPAycUwAEnzm0jKsYZ1CzSyk0x/x2OLmIvjbPJz7PewLCLxUFWZkdQsOPMGDAwyo2JGbM
3S0ENAaA7qXGMZ9fL/mcNqqPzzhPY+RHnjLGTliQO1MRvBYca4D950F3x1hmOQbBQJF7dfLo9ksA
SAAfY6v2ZGM9wqrGWC95q08nw6pXOl9NTQWUmq2SYIGB44glWfSDBp/1kkFW8i16ceUvuEE+TC+h
EgtgckO29b5IT81pUyZG4sadgRDdrC7NN8rcevUWwNpKFaw6bCwB3w/Ejr2FvEe6ZAPKn4zEmXjX
vOEmFYNxSw6aZyxm0k2kUZBrTV1tH0zs8dCKQT5NJi1A8I0itIn/9mCMe+xSZlO3cQ5amMZL01sW
bAc7BR6PCNrCQC2XwIIAPWYoJYAq5pj7XHf8VJ4h34mdJ7qRl9FFlfswVggjawgxvvV2AcMFY7s7
0p0AjY+bTw7TlwRAPKXm74EYBnPksNdUBTTWboHsQSN8PCwtTJzi5PY5RGfqGKA9VNcLn3pOb50u
0kFbeyvqHtLqShea+z9JeedtqAXMxwNyi+XzUjqgxrW+bwdE6WhJVO34aDqCQcgpB1u6T9WwD9Jz
9NQwPAYRRVY6/QhEvNy7jo7N6Tm2ofICvrY8stw9SP3OlT5s0d+NH2y6xCAt9lSjYJEvTEgGgvaJ
HZLnluxtgmgZuefBNNjZY1Uqjh+mNK4Nm/vMdn2vjurnlBW1/k5YBI1RS3B8+6BId3WZD52pQ5IP
zdcYvBQMcYsDU+GpygiOi8vAbsD4ddkU3/Z9o65BHa0WUcbgoSBiuuKIM70dTir/bljovbSFsM88
9I7u4cUpVutKi8ef9kaI+6NYh24xG7UwG0X7t5Pfv7TIZ5HYUINgxW/7nV7GJ/KJyuABgRYXRFm/
+KCoTbGxaWz5Bp92sYYi+7s5GA3inaIMpeKqpz/e+JilTgm4yqIHjcsNA86+Gsqp94y7qALEuvkG
XEZUETeV9rh1Fy8CItWG32/4tbNzqfaIRSuzBfSwp+kVw2h2VYO3IDFeX93JYl5Vdk6LZHVLNE4U
keter1Gs5RL6ILs/+iR3fVkWhW0zE/+YsQyPwAx7zTb/XmOY8J4u7ESN3SKaDL6FBpO4n16+yFG5
3A/Z51+aTGxMKRjJct7ABiyJxjLP/EsvcFucPKyhhlXGRfc11KaZ2RmCII3Px5JqnAWxhCFyyvPV
U3hz29DHvpb5QzNu2A5AxezTj52HTDqEu+JUaUd2t9IjbatQaG9PteOMeHQa0iTxwaEh1Uh7o0xn
q0bCxHzZ2RC4fR3TmFRU2ELLIX073h4twkn0fWQ/Hk9lTOuXtCMn4dw9PSa8IgbZWZR0/UgrbSvj
PLIBEVreTKg+PCJ3pZCQ8Y7kE1OZO1BH9lVsPetWyqW7l3J592i2EAjXGvfF7F2tA6mUwSHQ7lYr
4pwY/RDGdaNVRs3/067O88W2v+NHDg7ZyL5wVchqPZUiNI1FTjl1WD33Z+hbyDWAaNha1SVt9UZg
79D4KmehTM7fLqeBhsgUea3oC02S4+jQvcZdA3AMRhklDMC5QAbmWdZokovO53XImEST6S5DVYy4
oR5+c+8AOvXGY/1ku0nVFSh6VNV/AK+90eTaZgNubgwBPo0QJ1lV2kZU5JdPdkQqvPyO0H59dH7K
JwrrLlTFERTE/7cOhDCe8PopjxHU3WvulhHxUIgJAWIWjtOQP4poCp07IbWwvW5A4DIuvV5ypvTg
0PDGknkjrpcqDoyDRTVUVhI+QERxOxCPrUuqB15QRTc6NhmZcscN4cSMbO3z55eU6P8TObgo0/zp
ATNfRyMxdjihle4/1LT+BxwERsdlm98esZFRIBrEzx/vfISI3+mc6+PIbl3R3OuIkb7xN8BRl+jt
g9w3GZGzQ3gBeq7Bq+l+tVOkArOHN3uF84cLJZInQKFUqbnO7hiDG64iyatS5TIKsPLrgqkftMSI
eCdmrhhya5NNnZPr9tPEaUpnm5TyMT7locUlCzsS84+pFzNOcjFStmvMZkuY4bVSzCYGTFDdeuR8
g97sFeAoHzyuS9nFXrDDyn8Ifh0e/exQHX8lX6U2rADwVyC4E8MNlWgIzjdDlDr+DQGSyq8MQqH3
I5QfRJicb8inzQ4zpbimpLFOBgCL87g3H9EbF8vimlFu4MlLbW8W1iEbDfvI88wSprHNnisYnSox
OuBs2zkagelAUR9lmLUbsFGar6uLhL4EimydRiONpnhKs82XvBWNd6sF7+ndMtaA3sizXvtw2vW/
W62B+/GnUH00SZ78q3MTRfvTbaIZPJDftz0qY4TpkGhlRQ26aSItLVST1qUvblT1SvpPpOR5F5qA
xv3mIptMs0IdN+JNoyH9TOGXHOJg9U+G8GkLJrQXtN6ygDu6gXeTo0pM4sbIe+S0IHwBC/rZYgac
nhysrD9wZKm7gMUue+PxlXkJRwWez5rmkXt33V0S6S6iEtD5UEDwXuz3vOdq0t7MmyklIA0Sab06
tfEpHZXUDt6+SSVcLl2KERn4ZJvN8Tqdv3xdBrqfzP3Dq8cb4/F2kIcFqt6+KY9ZYZCTdjKmEPeW
GWv4wvNXfBYHA2SugruhDLitYWe2v61Nk+GEtsvMQz59QqXwhNLRY96XrB9sQ7Eqqko3p1jjRlAh
5e8qd1yzvZEkEuntzTHkc5E8TF8er63jNUhjIVV/pC8ytHWQMdO8cP0+4OSLmK9SyhwFisF08WKd
KMY0oFE5O6dZanXPXiKoMf+vslgyMQC6H4Gyspl7ufCGQkZOglYm3Gc6b/YkImUkvvLW2TsR2xSO
bvWToIQZvVkKYKURyFD7U8iZDrwepU8gcz9DmL3tnRBftjHFjPMt0ZExWc4nfA0RajwBVfKQRqaF
B6L7+kQAxkTtutn8rY1Zq95Eet7C7HHX0F6JzhSnQCjj3kfnkOacZ8PqXxXVfErdHRpzG/q2vnBE
L+Zn7dJgl5Z9m++o7w5+s5lt9AhdrGZjv5LwY1kzCdMOzAnCcqZgRdeOm40nbXzoA1Pu7OobVkKm
gVACSCZ5Vg5fBi0uzimcIjB7TxRFhRDU6jBv7rFzHpYpXhouRRJhMjR830mgRlPtEczmL6qW/odY
uawePz8RGVkjqSd3RJwOyLTXR36tnDOHTk3cA5nEW53BgBlMTlzQvLoz0FlRzBlYoQY522NrSCVz
kAQpu2ieqaCqKerNMdPuucwmaHCyX1Pgp9ynWIAtR8pJZXmOk7lAqEmxID3bQ83W2Ud9hs3iLr5S
ooN/eCbSV+WLAUB8VsIQkit+cpWzigIASVJr+KpNysodM/e1v3Fyblo80c8IjQ8EoYzwEIJV0BeG
aRhMXjVU/OHlT8sJMHBG6EvdHSTOmRBL+qWrZOcIjqxlyUBT41AQhwHUoH8HNm3cT0xQri1zgyUY
uzL8rIuaxw432gLDZ+pbjF53OqzSub/y04j4V+fXF0OcHKF+r/z3FZr7TbBVamSuA3H9WzWpJ1iv
LE8c/VWrbTecp3G4lwtYJPjFUzeG36/9wreEMOtRUzEzZrnyWS8zR3IrOwPY1NUPRIyld9sGDww6
3Nfma2gMOdPJyGHYcfG98kRhJ746SeUihOsW5cmxUPOnnblpnW1R1+VvDsNYtfHQMj4nTBna+HLJ
wQOp6wzibC83eiwJKOcqRhHEKu/yiv4v7555U2j9iDzUq64iwQsSVbRHJmwb3BennXjuE/rl+XI2
LXDmpbnk3oiQMXbz0GpHclnM9aG9ViMLDxgx80EW5a5HHKzI+ShWTZzFDhRTVN71nYyXrLQBlagv
XdtBhMS3Fu6OraO3zGbBZGV4X5BlQtoQgCZDbk4dQdX42dwLYWm9xjc8ftPz+28Gt/gf/5kCntU9
SkIGe/ubsoTa8ZqtnhG3F6cVyhr1CiepKb1a7hYNbm7xWbm/SDhEhQ5PdrEo+UT4EfHbDwR6XNud
aSEPPgK2u0JwBtA1CxmPqp3kcP2XJ3I5u0aM4iBSGvXmx9tZsqobJtqcNN4dhWxOoaHtKDlQ5XIa
tsrvMWBi86Qoj5q9s4nlm+geIHNYuWIglT3mitYGdOEqW4dDQOs6vyK2a8/D481Breul42JMiBpw
e4kO3JDYpQU/qBDinCFJlK+cD8kvQz9WZ6wts31BtZmQlJbvGOKcqmywXOsa3fLk4Dis7ydOSckP
MvfRlaG4yc639z9MyV5jP0l1t7VRKoC8qGiT6ccgeS4mC6V+ssWF+qP8XizjvmuZjCByQP8ZJkLm
syetZIs+Nl4WQSEM39rXXUWxFBU1CRtwsOchvK5q5UMEtjQxwlh54khE+/ewsB4CQ4ceXlWBPxz/
mULL6fbOIYtToeSJz1z627QMzjq3jk6wV9ATDH8A4ZTB5QEZFOfVjK2HfrUGWDSTwbYMf06DrUCG
ytWjQLZtsyn62eE4K9Ajnal8TJknMXjMFBonrdfhoslM7iL+2Ak6QsFcGPjgAv/+qd0G42CNDTiP
5DYQOPh39PMdXyLPpNR0stH291Cht2HFkbn5HHgqisQp3i7sGfmV0egwSENQNfFqAd6jZb5MNF9S
E9x4Eu67gXyeyvHwXOBqagIHdnfaxN18NwO4KCN7JEE01fpSy/4GmZK+hgASOwe8RxZPWbq1Ad0S
ISoDNOXx53W14vzTsRpxaJhatF5fI+jEnF+E4C0EPsCxmMZUspsmahQ94uvMqgNxm9WChHrHjjMj
LmP+Haj6djhzSMi7W5jxxlMIXGxKIxtUwAAk3gLqQmr6OMRzZoVU6s3gBfnszs5aBp/UJJYxParW
QpQ7f6zLybMbx9utugsG5Il7ZZj68q+w07VKwr0+I6NAi9ZP/YW0otD0LWWOYhur9y3TliS6vlU8
QkrhH/Gusxymjnry9IZZ3RNJdeOypYhv1cc8DmdgO1/4op6I4Oml3XoQqkBlqVFvhnGyMUo7XYgk
5dvCxm0uUUuCzG70JPj+kEszi0L2Q22wU66APuI1yDEdIrazCeIxsiCdeisF/pJOa/O6snqdsrUx
eUGgsaZ3wduwfPC9hV7aOhkvjc6ohDuV6JEqR65sfkuFtWmjCFJzHOajzuV8jJSgF/Q2uNVv6PAF
5/UB09elEQ6zH5X0oqQyeyFRZAlwrfWlR6Q+KG8bWR/WotnO3Mrt7Wr7GULvMk7REhg7LLYzQKmb
ZDTlsQm28r0RXnur2cK0qhhwZBIzn3u+Xotp1bFpf9CczUWZOJwzdw0hPWtfb8Lq7FQczzs22t3w
7Vzgd0KoIXi58u+GIGtixbe5eKReMjwJUe+6Y57FALZISs4m2uQg28RGfmCPBpj6UhLSnbpZLfvb
QT7eOQwjEM7Zv3nvSRbOY+gnk0gDVFUTeccz/tBYGcCdXo6iIgWVuPVRRsCDwBUAfqtI6TO3wthQ
u/TTzkeJ50gsoYZlH34y4c+O9XqvJy8s9iuxRPIY+uvVhZ7kC1Kgigv5q/VGrHB/3YuVRZEl3ZkP
l4bChQ7yWh8UHoDrROYBkxCJviQ3sw5DzwcVkynGc1bFcbB24qwip1o6siHrJ2hmWGAuGIgKVbUW
vxqeYIccPuEsv/55KasMS5Ncnym0sBNhkEUt42JAGCNn91tCOcGmBCWdcFFicA0N1MPWDVH7wgbY
MA/Xa3rGWF5qj1HWPdIS5GCFw+zEiGZB+vIPDG7MRoEEDL1AZ/EKCkGyPIGdogxyXdJafdfmSKZs
yVcJH4FfNoE6ymIIj4MVMcOZBPl1VNUgns4Hmw3AKz6Vm3s6GtKgNe/MKX/7NJ/2sFyW+LwbA3EW
ZU004Lgj68H3BoNysQBh3/0gDi4/7rXjbo1wAaUoaj3pOdA5q1FRxz+5pu9jdI0GQoAqYf0wms3q
CsFH6UiTRXBIfFA6lxbi9oBkWCFj+NTgrrpmu5DI+NPmdebzDBShPgASdpGO6+6Q4c2wiahQL+pK
VmskkJOM1rlddNbmsoJU4fxTMA0Yvjla48kIdGE5qQ68M8T3ejaACIzqsWEmw1L6LRP3UrkgHDG0
ZiIl0NjItSK9DV73ai9lr0NFPxEa578RlrhbzC41Vk32Kc17M+uFat84I/mZvcvc9l5jaAMQ9ELG
gL51o63zektB+iApoe3gvD9yTWy3VEguEYgEQ4W/PUxoJ1R33R9hb94ogo9pYrEk/APC8lqBW9GE
l/rUkxM4QGDya0KlgLsWFsSXSs7hPzuewlUARLFo/V7kzFfX2/V448QaJrNU4rg9M0KS1ECkNVzK
D6RHw887+qRaFczVDmQFhaicDKt33NjNyWEbTzKTH1rpMaWRhj19LA1XdpoiMCZid7A1ZT93gbyi
7UsezEHqixkj+u40QPXxb4qLNL4J16suZeyWuYFBUI9TMOT0Qqc+xSeW4O0ma50IiLu7+JhY7tEe
+Qw8VVCCcU9HbaMswmIsJRuQYsFMRQ1w8uD4t8cTlVsDYh36JIx9ew2+m58ZrCeIWeTO/mK1mLC7
4r71j/MAut8JJxYYZ5E9UsFYAP3S7mwJVvmdAV4t/KpykZhbfy+9+lnuicKIXdYOfZSJoP0+1Bol
okGF+6uNop3nHMjqqYds3DuxQ4T11Qk5Sonf4zCpNT95WXRuYr0xbCf4Wf/s4a8qrAdOiR3a2YQ6
TqlLjZk4wPOMQ5ARXe0Qiy9JHBqgo3O9TWzfwZ1fG3vFOKIpN/1tpvL9qEpOF0Jon21Nm0b2B7nQ
59pfaVC6cr61IV7Mpdk9OGIr7AAGENdxq6QQVscg8Nxpp3OJhtkw2xCe6fJ5BZSjkNS+sq725Oms
aK00Sxq2jRCv2Dt5p5/gRj51Whz03t9CBUAE2my0sQtJGVs83PBvkmAawwb8xC70SJEbSV3C06Cw
WILFhUNsAnh5r9pBxZ/tmMe5aT+MmEyuV0yENTt/xi6TFp1+5KfWQlIKgW5ah+KgWB6Z0DNATQyP
NssM4rDjT2NuQPRcezB7bCyipMwlwDTDyQHvbrpP8tkcewgHpVEISnqLWExBOVMS85OgeTRp0Crv
Ql1cODBtTd1OBpQMpqy7JCrk6PUY97aLEsY5Zzr/7YGmxJgSkFKvkuR5R0qEIBxANn0H7oSQWjq/
MYJDJ9Xphart1ngiVt+18OoCZYBkTVbXDj0JOvY2BUgz6Z4cASiVS3fzgZj3c/3HSdjMfPA5aMKk
WHhBpMHzrhxmMb2NCnDi9kPUvFWXVoc8zFrOZv92XNg+T+PwzEl5D0sti+ZWed5iv9jDHWd4Fw0W
ZgSWgRh72XRZmWbvOEtTxAtb+owzM+zRPcYi1D4bTAM95VzIan441qlQW8CIYskA4KB4nTh8/SIs
NiFkUYCltQerK+5efDRqAc7b/T5dXyY5yCd7gYI4ErM4RenY0uKuId005ChmGdZS2x/YmOuwsd1j
ER/PNZCcpV/QCmvoVoDiv5qDAbLPoTErMnGbMVsjQz6YLLRNyGtMrVu/XyqG2svcPUx4AFQ+sMq8
Zqkc+VtmqLJTc4bMVNIdd+SkbgCGF8caFY+YwlWFgXAEDjNkx6T+ik8Nn95dFH1LF8qajWaGJrOe
aStRQAcVuJmpw6aBcJVfb1mbUN4rsZ29TIZs6nN0hlGmTE3EBQqfk1v63AFjZhJ+kJSF4Jkbh9WQ
0wW2JALmai3dqyQpivv0R4HSQki+KBZ6fqQ2JsYK6TOxCGwFR6AoFQBT//NvhZvy+fCstzXvCsqm
/aOY+OnupIkboRRXX3ZOBjWg4ntdkmAVgBmzMj46rxnZ4ZcKaOeJwsc5vNh2pAs64fVco+W91EEv
5aOAB57eo0uwbtmpeB4xqNJvCenvU1a+ocJOM7CqABwYkdX8d+Lss1HEsNnPPkz4ysUY06opLvga
H0tNuVzE6497i2HfARBHs89QrKQJj6KRWuNRmzkOS+URqBQJd6HyQqdv8xiMW/9WbI+jwLI3wUTu
DcGHES1RMhOGFGyZnDuTpktC7rMcKYUAPX09iAvn8/pYA2ogZdICKDPCy7kjP3afu+uAofP+u+iY
KE7TTL5Ug528T3ys4kbHuHHqqOdY+nY9PXYIQRqe6GuSqsLDjiMJIdMJQjPeHVzBuWc+25GP3cbw
hBIOJhn/VgrexsmXzxUeb6+mXWQQZRLQXcHKKSlmrhcHQ8zYyGyTnauxmSboBrembhiY+ZKy8pNR
CGT3sjfbbNJJ23egFiS1tUVQQKINxtDu5+TtO2+vQuTWPaScYLyfPZGX2eco/dJbiPy/vUy2QwyD
4x37MhO3DjMjL6gjwYtCJ7ynqvAQocEvmuxJbgVisl04/fq6oaWXoMF1Sw0JGguFiCAX4XPovvOh
OUFBAhSgxAu5ajHAQXt8xrLI4dcDLek56COFUhskuavfmE1AokDqIlFA8p5kE+TY6DgX22R10PN8
hkaOkvuUqDqC2E+Yu0nCzLLWjOzg4M0di1LkpqLqQbhWkn10DpRg9/919nSYazKzZZNehXXw/Qg8
BTRf773WT5tCGInHN2zareftdVu3fnO7JoMSGsNkwR7WkexeJh662+RSD9TrY32YLCMjkQXssebm
C1Ma7ZKWR6Pebcs3ZNFmYQdPXhXBDgA9muirJx3INhs1HKSdU+uyGfbeLWIdyeXMwyliCdlVqG43
kWpTOibFPxPVqcY5WpixP1kAA7BDXnaelf3JF0mbZPq5qIkswtRPyzTzBZyc7pn9eDKl3NCi1NMH
VkPvrrR+DAi03EFY8qPuMTsBvebUobrB7ZKYhDH3r2Z5g7OgjDOhvp3ymqa1mrJyTAE0Z443ihYe
GstdhX9fR/FXBLiJQgRyJMaU56gMif8msRhcZVOPjg0GOOyya0AajO4hoDo5XEUtpE742lboGOPl
ugN/YkCJNbo+MKL0DUVNexw/lBoTEPa0eICKypGGl1SzjwI33ksQ1RNxDE1Yp0GDtnQWVUwQGdgO
+ozcRDoIw+PKUhpbWUjdr8zLwptdrTSkIlLAqS3rx9R4p5BUjLolh489mIWFQx0GMPmOqAkuaenL
JeC6WmixjHezHHiRGsLQz6VIZ7ieVZmTBb72XGMHHT0GMPrvgeIpnv8mEXx56PcVTZSl/D/R2UUm
xPVul2BvJ8wEzLB5FlRWRzuUP8kuMyJ2DcLAgQa+nTF64Fx04QzVAmMcPUwuvhFtBwz8Q6xlKXxt
0inp4GdEPCsGKradAHEesJJWflqmns++JK9rl9ge4s9AdVWxLxIlUmnFCmhVgY3ML/I163kBBrhX
0JBoNy3cishUNTaqnGMuM6zIOZ8RGciIj5RpM00yHqt6WL8c5HeLq5KwjnfSr2OrYlyatWfP70BQ
pCFb3JIeZnJjCBJeQa+49rDfUAD7Y6MESumKPQejZkvFWELaiNq89kFTDbhjcxbr/d6AR8HXsEqA
++wsvbzpqW8dCSfkgX9pl3++VXRrzeFCzNrXhyKDsiTkgIGBoULI95b59QnUNxKNvptaS11aw5dI
XQLLP6lZQ8DCjfearkjuDAqJiy4//ONfhYVEQxbn4fzY/tx7P3EsRSkpyBMY5hj9dL+RjlrVRWKO
APjrRMGpxt8oNW1Qq/ejlWczQQB1ogMfH79rMuRnvwx29AK30XFToEGWggAS7DKVbwxHwC1+S0hF
8KEF9pm35uaBLUBwGvRrNUWgnoxP/snbVDkI20kBK1apL4Y0SDSv9JWSkEYTgPBTzgKaBRQO28sq
o2Dz7HwvXkhRWovurA3wsyr29P+pG/DV4ZgEX+gk72mYp0LavfM+0IEkQJJNCLsDZ62l5N3e1kqB
W1lQINuWIm+6GEcsTpEOfRWMl17dTRe3rgGk21cTV7kdqPLw9He3ETqvVC3qsQyZ+v3fvSJL+M5Q
1YgY/mdX2D0MM2yHUj9vAAWUznbxGcs7B7nxgIPg+Lhooziu5LYtNpq/TEehlZ+du/9DqgXqXoLA
vkCxYx+Uqm2Xef0jC9XbXh/XRggsp+ji/I19O379UtEbud5uXpvLoIL7IwXwjViPYZEzIBAm7vne
L5sD/+zPiGubtQ0nxWJudQhY3YRX3sKuwgrXlcS+3r/Tx02eOGORPRtZ6q/aqQB+2MWCY3vbePIu
/sASnS8G2PLw2xQEwD4MWBJ7i3wXD4HmM7P/TDmQA03pvtX6TJsLh6+/qML6Q0af3u5oLMUQPgO7
X1kffRodJM6jl8jr7FmiFONEi7W+Q5h3bB+rhlxNEM714B+TWSWvOva1C1V0UcitiFvZJQYY6kQy
biNivcI=
`protect end_protected
